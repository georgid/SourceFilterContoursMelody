BZh91AY&SY�4��߀rqg����ߠ����a�o���
�lA!LZ��
 : jiJ+ �=�1M��� YP
�5��� �s��QS��QE�      *��TR JETR� $m�̭�E��((ڀ��D������$�E%/&�
���������$�E"�H(�M�b
�*DE��`�R� �  q�^�Q (:�
4���.mva��R�n�4�]j�u��Y�d��)E��T���ٵ�̻�˭zuʁ�F  ��  �ot�4҅R`e4 �C�J6�ڶ��sT��F���@���Z@�s��U�C"�M��u(��vFU���c 	((�Aࠑ��Q� �� �M@��`pt	QY�UFa���a�T�:UJ��t� a�wW���	* A�'`2C��2������fTh`Zl��0 ;:P�j���x �@A�|> hf{8�Ez��\P��EM�(60�w0���@t����ڝ����| �  �p R���#ۧ ̱�h�
�S�2�);�{�Эu�
�iT�I�.�]�և�� )E(� ��P-b@�(
����s8$��QA4s��KN8A35R[6�5�@�6$ �Q@�E�0�:�M�������������4�ͮ	�v�A����.�C�1z�;�  <�t͋:p)ӎ�#�։��� �8�cn.�nۃ J@ i1��Ej���x �T)xkA�Eh׷B9LFƢ�l�4�`ѭm;w@:ón�H���                     �� R��<�M�@��   �~�R�!04�m#���U?�ߪL�T����4h�h��22i�LA��)%R�� !�  b` D�T&��U0` �0�  B��J��z?%<h�j4i���i�yL������M�������� �օJ��K6K���^V�P � {�?O���Q ?#�P��v
(�(������?��O�bï����_���0���~��_���������������;����~[����K���r� w�w�r������?]�� ��_�&2G���?T���W��@(��u�������g?��������P@@���S�I�=��������J��$Z��^��:��⧈���q��:SË��Z�O�#i����>�u󠱺�v���f�[B�*���F姮DE�wG.���������ۡ�jT����VF�4���T�k�����J�-d}$�0>����,<eTn�#�Q+{x�3Nm��'��&���� ����o8�����n�P�jT��[Rø孑ވ�Ȉ�e��嘏1�z��t8��VQ��*�,iɕ��J�2;;zR�t�@Fn<��'��|7f�@f:��w�)bOl �P�`:Q{F�\C�R��y*�P���m��F��6&ro*�Ÿ/Oj��Q{�ʌ�g.�S�(�ܭ�!(�G�l\N�JV���l�ҏRb�N��Q�)��b�M�f�@��}�*��Wʲ��=ݷ��J܍g=�#��<+�Y,2�n[�,R�8��k%�-���D���7qlX�2�4mb�D��جղ�e��.�V�S�5��� �)�w�/��m �gUJe,d��Σ���!��C�HU!���z-��<ȳ�#�f�lV#�UU�0�(`R+���L���w�K;��;r���ܔ �Q�i,��wUf�!���~+eJx,K�1�3o3�����DΛ�=�E6��v���F���6��Z��Z,m��.�ij��nQ�W��u>�9�8e֫�CD�Ӧ�Rj��$��-��\vI#*���H��JWV�'��b}��vy���S̓Y+$q�5b�a����U�����(��U�1]�R����E�J2.=�U�N�w�'XY���^�*Y���v��*�2���`"l*�U
܋"�v�q���U�]ݴ/Z���2��v�
m̔3�WL�f�$�7#i��m��
�ҡ�:��;��Tg���p�e�f���VVK4$��j�P���(�扮�j���]g[�y�r{���
�;����C��Y!˒Hd�d�w�5u!퐞�	��9�'��s0n�:�*�H�а��܎ݛ��hJn�zra�Ô�7x�y6� �Q��/�:r�@�X�k
�������{�<�mS������5��V��x+t��vs�tu
���S�MJjSR�JR��)Jy:��kκݬz���o~�'t�n�i��-p��y��E��k���u��RV�����-	��q]���B���t��:�c�9H��u�{��':��ڤ���)Z"�P.�Ʋ�w,���^\LG=�>l�N�#��C�h�9� �����v&�xyKG��"]��|�{�_;������G�����z�R��M����n˫�dj��7�}9�|��L�EdoÚ��'��{�cR��C\�g��%��%^c}.U|��+tuz��5�>��w�|���5eV�F�K凑3#r�P瓽����1+|�{gG�c���"�S��}k3�Ùg���r�yN�t�U\��c�>�[�]�E�y�|��\�~�չ���\��/y詉���[�Rv��Z1�*r�ك�iy^  Bf@ )�U)ݨVJY(wd��JJ",bBf�K$�ڒ�c��E=X��+�Y���G��,y=���F���v�ְg~�F��3g�V�}^o�3N��)Y����c��8v���<��յ�9�F.���+c뷔^&�����u�yMy�vv�ι�k�v���ce&ڡ�R�/'&z��%�=2  ��� ��f@   �� �U  L� 
w@Z�9u+�w����̣b��E��_#�V�;�%N�>U�K�u���;��b��G��ǡ/%�a.���fnNr��[��}��4}ʞބ, y	(^�lt�SY�U�My��37��1+Y�U��Z�Q�k�{�z�1Ij��}]�)�2�l�V9��:/S�;�)LvbgnY4�h	��%){.�JGZ�UR������)3�X�-"�]F���r�c�TLϛTD�Y��3.��ԥ����g�����5,S�w��J_:���Mr,c�#�iS����-�M���.���ǥ-��(�|�^����N(Ss]K}u�%�W��9��$ �C��H�l!����FNb@��cr1(�]R�c]�u4MW[3��H;V�ׇ��n�lF��L��R	xޝ�vU�eR�l5��ve%GS8��ܬ��)eC�Rآ^�o=p�(�n�k-ʸ���)/t��P��jm��N=�ۊ�OI�zAJ*ܶ��J�UE�ʄS%M���Ǡ�p���J��W�A�U5��$�wu&^���6��t��apKA����mѳ��)�1�R6�����#�
"����t��)Ec@Q�b�yG����%LiWF���sF#��C�-�9q#�/lc���E�;�r���f{^ڗ{��p�S�JK��
S�*K�H"%�rR�9Uj�D���R���'ϖe%�Fy�u�X�_)�L����}n�1�ŏ��&Z�+�T�d�V��K9�G�%�[��l��{�Ž��)���j����/�5-�ऺ��|�'���[��N�1�>su>�:Ʃ�ߓB�<1.}�|�<ĸFC�����1�����c_:��O�k\ǄG�.k댖O5�䥫��%����f5�X>RrY7k䥇��N
<p�6��U�p�q� x ��m�Hp���:�|�&/�R��$�Eg�����5�{�T�-vN��3 8Y��(�M�Vi)k�9;���sr�w��;�2�( @�Ӿs�n������O�2�5�k��Iԥ,;-u�ܖ��
�G��
6�>^�L0}(*>��֬^D�|�%o�%[�vz)My^�������O��^U��Q蟝u�^���,r^JEd��y)x}�����ĵ-|Ǻ�'�k+D�I���y�� :�H���)��[���)Y�3��#�8 uьr����8ɜ��{'s$ɢ�|��ua�s�0�ZQ�i�ģD�j��fu��ǸYEh���wU�f����P ��.��������&I]����J��ߞ�|�mk#y��  �� �À<>p��$(��R��J#��vh��f�`�%����8�%o�8˵����D���q�J��LUk�s즫c��;Es1�뛔ş"�+5�����OhO=�^M����-��L�]|��lM0ݿ����(�_8�|��)�Dӯ�W�w��b{������r|�E�O�z&Z�My*TVD��X3���W��k�>�q4��>S�,ք�m�ʺlف�=�F_0�p+=����J\k��&�zo���y�WNL�=U�4@X�B
� r 0�M�vZ�|�!�m�����(�\M.1M`vQ�.�c��[k���Z�Ԓ�^�i%D}U�}Mk�6�=澻uM����u��מ�:�'z�<���V�j��^lnLvyޟ)ʜe���c�n�^�_>J�%�L��2�iT���~S()�Y�3��y���op�:p��,���)�UډE\�5mS�]DҘ�9�D����h�(�
��w9��#�ԥ鴥�fn���1�^w����r��Q��ui�51����c�$���2=Q�Fvu.��J����樂|����	6}sԩm�c��W�WV�;�R+�ՋE���|�1��T�L{mb��:��M����k'k�J"ζ�iMky�/�X��JW|���ϔ��.|�1"�l[�i<���:����u�8R��OD�m�_{�2��RR���bV_�w���K�"�ǆ&��&-3=J{u��ui^y���D��u��}�G.*<�=;�8��eN�z���A�ޮ�d��8Q�9��,��I��s�Ȟ��wK+w�S8Fj!�%�h-ێ�]׏N�S���R���Sk6�z0Գ�F՝�l�n:b��X���.���wz�x��Dۮu���[Ǥ�����=��$r�i�ΥIb���%)ɏ;n�W)|��R�SnZ?5O��� ���y@���>�-�T
M���Jk��=��|�%��m�Dj%�s�ח�>|���y�߲�)J�b���)j[Q>S���OL�"�$��g��P�l�Ed��tK��M9��Y��M5�u��y�5)y��q2�S�����D]�jw�E5֭�G�T���,�6~��Fyb�)鉎�O��%.��T��5+�=P�:��)��ʱn`�Z�ٷ5Mb��lƭK��LP�#����j�kF�,d�"�Auçw�/��,�� ;P���P���5�M�H��"���VƱK��c�u�Z�w:=�AP*}MK�����U�X 	]]X��`>��(�LHc�#�`��WuBR��)�b@)�#�u ��,Lą	r#&yrj�J�v����T�ż�"PK*؋�ΐ�c�O�Yߔ��v|����I���(�Wf�מ��,�Ɗ! j!G
:D��:r�G]��V��+�0��`SR��P��m;�n�4z�n��*�fZ�e�'Q�!V��K��G]����2��ѝ�u�Rc @FT9��^��w�g[�Yl#Ƭ�D?�U��eҸl�����T�k���j�\���ʸ�f|�$_Qs�IV���.��s���E�?Ug���&
����j��t����S�9Gfc00� �wz ε<�s��ܡ풇u(wd���Ab�⸉v9�,:"��^���+�v�W)R��0��Tө{����_m��Mb���o~s�-�X���}�1�{:ʋ�Z�W<��/��Js�w��a�2�ĥ)L*������M���.j��I)P��JR�
J:�ͥ�%JJnffT��"I��) sw6��3*��X�").r#Q���Jd	��2�Uʫ[րJR��Z@���P���]�bD�]�`��^��-)JG��-)JR��ե �I^���gj��H��ɞ��ɪ�ى��uxc��ٕ����K^�UV�6�P�oQ�L�d�	ܴ�<9�Fu���/�!�P�����$-ڵ*�H�f�\W�Sic��0>����<��{т��-�rPx�Z�l�J��O�Zv�0�6J��5����"�0T���>XnU:X��Y�&����8��X���p�ёy�W�m���9��휕�"a3��|�'EP�%N��^Ωa�{�a�c���ɂZ��S=u��I�ac;)�?@���i�ݔkOi�m��kb�oE�xm%�x7V��c���E�.].X3���(�}�1��>D�"3:HqA���0��\���難6�\͛*Sr�RR���?������UV�	b��b��nn ^��fC���`�$��#��SZg0���雃��L��x&�i7b��mc�%ef�HRx�)˩��<M��LJ�f�����=��)#�J�.�8�w��H惾)�/H��(kd�Ζ����Yߦ�7��Y�J7��O�+ħ�tB{��	��:�Y�s0ߜ������"N^����ch8���y,C8�l�ț�r���0lͺ���߷-1��5�Lg�S�n\�V�;/;F�0@�����$]qEc�pz��b8�dsk�rފ�����E�}/��:���XժǮ\�����zxWm^7������])����[G�z�T�?���>	u56fV���F�RZ����<�lrM;�Q��WR�vh�#J�^�qKɻ`�˺NI���Fpg]��w*C~#�;B�t��"��t�\�LQl�1`�K���vj�t���I�����ҕ�Mp��%BQ�}�t5wԳ�p�A����gY�䨕����q�b�}��7\	-�%k��1��wq�b����r`����]=b�B�D���D}Qp�t�4j�U����n��<��V�+��Rи��Ts�����
um@(�U�iWj�dSqR��&��l��V�ȡ�Z��kw՗0ѫ���<�g*�X����Cp��5,]B�v>P��q�
�����J�avl�������Gk��@�����U+�����b}�����s���h��bm��E9T��t^��!��L9#{{�g�ƫ-f�X������uE�I��˦�=꯽�ݜ�E�5���/L����̬���223�����ddw+��z�Z2222222222222222d��U=w=#��FFC�}����$��VJ�෽�� 2�]�o�����2/#b�w��ֲ)�����FFEd���dddoё�{�ح��\s###~�����bo��y�܌��zdd��%�#>���d���6^�#%�KFF}��^�����輗Q�v��M���V��]�����v�qk����/�v���ܝ�ɖʏl��ww�絚�ϣ###쌌��ffO����g��7̏�22K޲2/%�dd�%dd������Oi�9�jZ[��T�5�����_"��n>����w�ђ�/'�N���Ƚۨ�˗��7}d���d����d���d����222|��ɗ��ȷ��*K��{�h��=�3�Z�_k�|�w���c######'{�Fr������k#########&쑻�$mܮ����FFFFFFFFFFFFFL�F3�M�##=/���Gr[$�n�_k�����k������r�L霠��WF���[է^�� [L�e���㺍5QꢗK���*�E�6����a�m�'wq�'b��ǆj��)2N��a��o7z���2�wN$�3��ۼ.ʹ�rK��|�Q6_���=�������+Vj�gbZ������҉�|&IS/R�������r�zY�x�[��8�7���������]��s�n��on)��]��q/zo��3wJĻ�U���a=�^�)���ڑ�/��m�[���qY���p��ގ�ow�mH����XL�T�=�-~�ߙ��M�n���]��2����ww�I�w�� �3;=���� �@  n��W       /w`    .���  ��     [�W~���m�I�@s*���8Ӡ8(�̐z���뻻���N��X%�݂]ڪI5�} 
qrI.��I#�@pP ���r����wvS�ww`   �wv  ��      UU   $�   2��� 3;��<       ����  =�I/w7e��%�݂]��%�݂_n�/2�U}TUU���%�݌̛.��9wv���K����$Â�{їw�ؒHm�݃o%o  ����뻻���K������	ww`�wv����$�
��� ��S����v���e�݂]��%�݄�} �/2K���I�{����%�݂]��I!N�$�I'c�8(\��w}�υ�� ������K��$�z��ޒUU@  ww`ۻ����8Ӡ8(��wv
p�@�{$�K�����K�����\ۻ�]�w����G�$���     �����   �$�      d�   ;���       UU     �  $�        ��ݘ         7w` K�� ����I=wwv	ww`�w ��z>�@    ��    $���&���I2N��> fH�wp=$������ww`�wv	wwa.�� ��9u�/��{r�p�8�{ي|�����Rk��P��)]N��H��,��wb�&v��7�I��Kbl]+1��X����+��ys�'wٖ�����׻���;.O���F�J�z7��j���&:0�6�� �w}ܘ���wV�K;���}�6S�Wh�/��O�&/{�h�t��}�m鎶���lƪ����S ���5���5�D�K�5!V�J{N�;�%X�5H.��s�"f���C�f��Z=秶�X�SA�h�x��%�,� �Z����0Pֺ��s�ۼwaPb'Y#��ր#t��o��-��3&��qa�8�N�&Z�օ��ZN��%y�y���9l�Ac��I��eґYGZh%��Ų�/&P�$�: �YB�w��-�;ZL�Q�*���TQO7��S�r�'�ø�nes�6�U˖Wt���`�eM���A�hF���JV� �Kܾ�f��)V	�uu�Dέ�cA�MoOQ��^A���F`�:��޻�EV���@з.j�-ګ��a�j��5rFչYR�Ka�M��"�k�(� �)�&$l�KK7B��^e�GL���̨��{y�U�%Z�}�T�_;�����V�UV�t��mc�ϙ��M�*�r�(���:��i^*���O=��j����[���ko �U���3�7�I]b�&s
�Y�vTXb˱ZN�T�0�n
�'-���"R�6�R�tn�gC�ZUtz�cT&�uL�k���3����0E�(�,�� ��|v*}O-d��5��~Ssr�q��o1�;ts�r:�����x��kz4����%Y�Dl��qۡϦ^�ݮ�Z�u�	kTdp�*��Wv�$�ܐ���U�t8�^��;[Ӫ�ǣ���/k���0N����WF��G���͗:w	֟J��{d��ߤ�Eu��7b󷤈�#�-2f�(w���v�o�P��hD�yliە����l;2h�gX�b���q���g*��u���f�3j�d�����e��-��vcaV�>��4�8��%H�(y�M���+a>�1+��],��+����$(+��P�޵��.���iG�^eˠ�7�цV������m^��jT�n��f:�h�Ԡ���Q�t��&WV��wnPO�k.�u����m�;:��|��w`ߠ���c��:ng���P�4�a���GPS���b�Q��9�o��kT�ѓN�Vz��4��.��J�[9�ؐ#��(��3vu�[�*{���y�NZ���*>�5Җ�$e�S7�W�Lܒ�-Xx�5���p#��1��n_u�w����&����i����Ɗ�B*�mH[p��@�S`����h���7	�{�.��>���n����XoSs���7n��oD�]���Zu�ʤ�n�s�[�"��f�*�+��G+!����7�N3Z�]Чy+;����꘢�-4�����^+��m�(l&켶���g�Јfʡ��3��δ��+���m��E�*�x�ݷ���7'��hֹf�76�'�=XjeY�L��F��rd�֚&�`�\F�z}��U-o�W�k�6-R/.�e���2�%f��ηY0�T�e�b�	2T�eؒ�2���1�^싺m����:���zz��#��9��9R)$
f�N�E'D����r�)�d*BpH�y��n�rF�0༽���9-�q�&��������n.��ڼz�����Y�&FFFFFFFFFFM�#wvH�O��]z��������m#}+�{&�%��ː�fƁ6�o[m��k�9���	C7���(���S��[=�k�x�z]��ܛ�$��ّMWw5�;��'.�m5��܅�����*N�ĕ�t�^�V��9�R�w.B��Bwb0T�rk��E��/q��(e�ۻ�wt�g�ԡ����[=�O�۶�r�+=�i�&���fG��z�8x���EJ%fc�ծG����Ǥ���X�s|�(����\C6BI'^(�*4����Iۮ%JI�����p���F�-�38.뉬������z9�^�z���W�ɒ^�o{|��n�22|���ɗ	su0���׍����#��#�y��;R���J��;r�co_k���_k�g����KJ���_k� �t�9�fE5My�{{�z������}܋����:�yږ��ɶ�ؖˣۖ�W���꬞��p�d�ҥn=��,�,e�WoH�.��Ȝ�Jv���}r�z˧�Q]i&���eYˁ17;d�fdv�KrM�i-�f�.��db��	���}X8�:��ݻ$0���FJ��)�����۪��3�6so����Ď�Z�
ǩl��_k��������ۼ4o�˻��"�wg_k��fɯ��_k�����6I5�q���������zA+���{=Y}�������{��ya���j��y:fL�3���2Ew�L�<w�N��j���˙g�q�P�2��׭��d1�qIjm����PI�tv�Vv)+3���[���X�t-����D9�H��b�4o�O��ǀ��m���r���^�T��r�����
����1�J#Rv�˝$�w7�fВ��K/+f�]Y�zg"j�ݧz�]�SgkV%������O���I$��nw1�fM������;�s��y�Ͷ�ȹ)w9��w�.�vf����Д����ov�K�3d�5���L����>��&dw,�I$���8p��_h�r��y����k���F�&�>��4�`�����|�5Oq7�c*��M����g��22222>��ۭ�}�[���[ɷ|I��Z���R>C6I3\}��{:$�l��`�b׮����V.222r�ok����c##&J��FFE��s2�u�{���םĹ�kul{��v=d����$�l/��$ًئ��u���i	p�I��v��k�}���w7�fE�I=�v����LsP��}��� I=��n�c����]�l���i%m%���P�ZIjFk���I'\�����������dc1���6���3�����̎���_k���̖��$�$�$I ��-Kd��L{Zsz���$���|5�F�9�o	q�P�K6�fN�]ֳ5���*��Ij��KR$�ڻY$����$h�v�Z�###"����ʼ�_�s3�ڪ����&slP�m�f6���pݔ��^���) �K���{̂���AE����`��H�v5�d�n��@��w�`�.�OWe�yge�����q��ɩ~+}�5����ȕ�+ޯ=�FMޓ'�wf6�fϾ��r��"�x��U�fX�yw��3�'�ffH�dv�}�k5����������22222222223�wk�����������U�d�7Y�1��w����O���m��&�22n���F�J��H�����������ȍ��EfU]׃#.����wzl�}�2���Q�$�%{UA:䫝,�-7����ٱR
kV�[wo`˨��;�
�l���v��n���\o���.x��}���]��V ��R���eM�ͦ�\$�X��6*F�����a�m�-:��˘fL�h'��5ٱz���Uc���EuM�`j���aXg��[`}i<خ+�+r-98�Jy�C0��L-�'�|���ZVVu������b�@�.j��O)��`�9X݋�	�h�X��>�C{s3E��k;��Ъ����E.�WT�׋;��7�"���Y�F�l��M�\�N՘�s4/�aamV0������u�����{6���C[�m��۶9u��h鏴�}�wQBl'o�� >z!j�t˽+�{�j6��n>��|���S�0��m�V��mj�oH�v���[���bm�=h+��X�njV��[� �]�;�(�s�Y83i���+�;Y2L��뢪%H��u޼�љ����v%sR�}�ܙo��^j��"+U)R������LT����crS��\��s],L�陘�,K�#Gc[bM��2�����������s�����V��\�!Gl�}�:JE�e�7Y��v�\$��q�z����ݝ3@.odUt�J�X.�ЋD��烫e������CJ�Kli��{N�U�a;"�<7v��/J�o4�A6m��C�.�~�N�w��0rn4-�;1����vr�%�U�[&���t��Emq
��lA������eV��r��w.����.v듇k�1@�ƭ֟Q���|�|��9���ޥ�b�Ȼ��.�����w:�^ŵ��vv#��p�˝��j�z�])�D#:�S��jv�r?���\�\������1�}2���9ueᝯ��Wu��bm]��Ά�r�T�5t��A��R�n�Nf�3"+$uJ�I����s�{�6z�tJe��V��RLk�䮶�����΀}�!;�0Mn2���.뇺߬�6��pY��r��Yc],�3;�jV�|�u� ���
R��Ք��8��y}ϋ1fm�i��؁��]�; ����K�'u��́1��Ȕ��Z�A���&����uȑJ_Rz��i^��{(��gʗ5�Y�KA-z�,[*Aveɓ)Lc��=ӡ4ܡ�Y�qLs�e��v�5�`8pjÖ7���I;�SҶ���'�Ūӻzdk)���*uq�����ɮ�����iι����Мv��V9o-0���N�63�<�P�yF�K�J<�����[�W�7�����ҽ}���XU�V��q�;d��v��O&_e�|G#&���ꫩ,3�g�X��|h-lݤO2��d0]鬝���Ƞ��G)"b�j�"Rx��V�
@���H�ʾ����T��R �A@�G=�u8$�)�-��x�-��8�_X�]�7w��pC.4��k��Y�}Nr�1c��	'�V�ސ�ǜf��9n�QX$�ё["�<�����=���	��j+j��*���#�K�Qw;h�N�i�[J��Y�#���^�y��o]�[N�F�b�ή�)υ����]Kn�9su	wu�W2��n!�h�]ʫWu�X�N����܆l�����[b�r2�Tv>e�r��}o���ֳ*�`���4Th�ƁZ���8v�e��v�җτ�^�S�z�w�]v��О}�c91�t���t��t��ͶξVM[��&b"K�Gir��.��[�+~��7���'�!�;��q�cd�v�in
��%��e�7o%��q�=T�x�T�e�A`��I�|P̹}�Վ�q�Y��V\�+z�'-ꛧ�GeW��������/�/��E�~����N����������g��9��~��#�������~����}����1F?���d��7=�r�&��X�s�fU&�v�zp�*}*�K�����#Z:�a^.�1���ge�ܷ�v��S#��]v�bx=�"<�z�@t��LT��xg,��ot�=z6?-��z4óv<K��x/y��m�S�q+��2{�f�'cz9�ۡ��b]k�ӎΩ��3�H��[[�ͬaY��{W��U���I���,��9��s�0����5*;Ki�J�H@�X�j4/��:�����z�0���yV��sV6S�f���Z�2��Y̋��sl��8)W�}U�>�'� ���\��ǝ�%TN�H����[>�ץ��<=�(� �/a���@k�j���s#�t7F;m�&Vl9���fz�$"7�S��{�:�P�X�+��L�S&�ч��$]l�׍�}�al��>z��6��Z/�C%o&�Eb̷{��BI�פ�����b��>�T���`�k�[�V8,��89��a"�bJ��}_<jPi�Y��Pcx�r��������8��{޹�qu:�<���C%Ѩ3��\�b�a3�v�r�p���q�ͤ�}�%�C�Z����WaD,-N��H�W����v���%��f�32��u_|��,�(��e��=�t��T!�_D�5��"��zv��>C�R��]]���cl^��ܒ~���:���M���|�K�3�x��u�$u�&ّ#UR�"]�V��,�(rG��a�j��Ll��H�5u�V�d�W�[X8Ύ��T�֎(��g|�=��Q2�4�2W%&�Q,��r����S9�(e��]�g���^-D�6�7-��&�RQ�هv{q�d'�C[3��7s:���
���(�F掬�nX�V^,GNS��HO2t���=g���.ǩWhk�n���^�F�ȣY³1�M��hFS9�fҽ�q���@�]I��oe��X�LһA��ç�.���9���.T^�"����,�u^9��^BVV�3� �p�h+���
&b*�R8h�&A��ϩ�3Άc��府8U�\F�ږ�g�wp��ܙ�:a�� ������Ψ���D�-�~�ּ��|`m��Z7��R�]7KR���}Hx���hkrGUܳ��A^�u��'"
@�E��N�u�sC,�{E2�����[ZZ��W� �j2�_w��YUU�AV�9^d{���v2�ft(�j��
�w8%T:�v�����������KLGow]f��v\���+���CN���c��)�8����Q:�\��ɪ6c5(�pP�|MS0W7����R��I� �;�vYMYwW���f�on��'[|S��3��Ԭ2�d����ųd�[WIV������BP�=�)�0�{b T�Y��遧j��sݧԽ<6���Տ^+�L�V�`|G�8�xxU��#J�nr��B�ܥSs�����vhvnE�n�V�oni:�Q��D_M�\gB͙
������ �U􂺱��^�$��!YDʠ�D��╚��:[F����v�5��2���o`�����k��1�| �Da�m�{��/���5�v��f��|��J7ٺ��X��y�K�|�V`�x�?�>T��N��j;{y)�Kx����Y�l���P��ʇ�"��+����6[^�8AMˋU4d�e�H���ʋ�xA #��y�xB=���iS���w3�*��XA\�sT�����ZW)]W�mN�}�=՜̽�
+��[�N,"G)ja�\�y���O=ѝ,!��j�������Uu�C�I�r��+�㯪�D�"1�ɢ��.��y8�2VC\,�t!����,Ύ�G�k�]�	�R#��ĬfsopL}̞��#��!�Z�7�-��ʨ4eM��ʰ�E:����`��SU�N��H��޷H����R�UN
%�.�c �hi3,�-uxk�SM�_��,G��]��������DI��шn��zs@�en;���Z�PGg4���
�߱�ɳ7n���1\�X�c�m(���6%��PL����Q�=RH���tdJ�
�vP����1���7��'����w�ԙYY��ު�<ں�����V%�u5d�yY�ȼ䖂f�Щ��������
�8�2�-��c\K����UU��_[�S�����mq���I��q���欩�J�/gKCebFVm����{�������r��Z�JW]Ѫ+�QR�Hևӊ�jű4e�YU'��P]bGtO��<�B�;�ۋ�u�\�<��'H��}_�[�n
�T��6��Y�LsR����4��uffƐ��+Ŧ�'Ŝ�tۈ�3yMN͡�_Riжd��$�'0+�K	"R	���vh���v�'�Wex�d{)���y2�N�)��y�O�&�������P�9���"�Z����6#�]iGpƻ��e�7߾�����
���b� Q�'�׌���yU�r�`��DUP�X�
���ڧ����6���!]w�Z%�xS��Co������4�K��D��N+��V3�m��NZ�,�\�*��Gܶ�L�W��QK͊r޺�z���I��r���6>lۡ#=�zd��\mmʎE� ��z'��v����|�D�Uˇ�πC`T��AҬU������z��l�]��W�Yr������q<�)GVl]��/�#�.:�uʈ_��oI]s����/2�|����q�E���ol�J�f��6°�V��5Ј��㵐�v*�	섁�.ї�l��-;&M�&&8���<ny�x�3l"oś�WL,��+- J"Z�X2Fe}���Hn�S����,�W������[���lt{)-J��F���жsW��+���"gm�F��#)��y���\dmo����e��)$	;@��=�}�2 ��U�2����S-ojniAwcÀ��� )e5��Dzc�9�CA�KZ�{6��V�/f$�wd�҃o�g+�%p�{����?n�1Vړ:��ߑNw�3��:xuj���Ǜ��3)vR��&۫���_jH���V�]=��[b:�2f����5a��d-lVr��^���w<�Ӫr<�¸�^�҉ W�3��і�h�J��F�
�C��^ F��ڽ��gh���ʨ��xY��(����A�%
�Yy����b���^�˰��K1L�5^n�����\g7�Z���ķ�Kc�9�]��|����ٜ�r�a�c�*;5�VGx� oq!��ao*�k���Y���!�2�v��+����;�)�e���gx 
�Z`=\  ����.��u!����\����Ú�n�W���H���{1`8< 9V�.���e]�W]� '���c�ѱ>�C�6^������	�~D;9Y�t���N�w*����́v�C5�������r.�Ta�}���J�O���:�5fr����bcm+J���lH*����9d�"�\��t�m?T��fԨ�gw����F��-�1�2e�V�N�:�%j&2�\%R���{Cd�ۗ��XU�T̸��J�};`Ǳ�Ww�	yIЭ��!�n�ݻT����#�S]n�-�|=�,�D���部0���jKV������Ǔ��o*L$���!ME����}�/iM�4���5���r(�;7M���GGJ��k2V��/�J�N���\γ퓣�X=�Vv&��#��\�cB5P�먒{t�+��O9K�u-���{	J������j������̓�n.��7Gouua"�oY71q���Wԍ\8֛���8c��w5P�A��RI�'B���)ׂ#���q���R;vowd��#i�$=4.H��k�[
EB7�𻼬cIPsR�޲�^�wp�x�G�MC����n�A$[Sy�ھ�Pr������z:�k��������� L��>�^��k�f~�b�oW�c�����R��*�b��)�h��������̨JR����U(JD�h�������   � B @G"��9�  @            ��U UTT�UU      ! Á@@D$�H���((������   B   !     @  �  @  �   �9�   �9��  @  �  @  �  q     B     B     B     B     �!     B     B  D��@B �̂P��@Ҕ�UUUUUD  � �  B     B   �  @  �  @  �           �  @  �  @  �  @  �  �   �  @  �  @  �  @  �   �    D��    3��0       �  ��             DGr#�            BȈ��  ! @ !   r�D@+�@YeUTH��r8r��  ���*�iJR��)JPH@|<��Y�2ӉA F�)$�8L@�'���H�^��$hG�6dl�ڑB�Q#&#EW�7�~l��T�UW> S��{۰�ڀ �d��6�����OUn�@e�{޹= 8���`� =� }��U�
�� ���zIw���;\��q��қǛ�\�I��I������A��v�f9�_��9H�Go��x5�ooe7;�g[��D��.���<�4��R��j�E�5��X7(�q40�j��TGn�I�ڵ�*��]�譓Y�B*o�T��>{�}�j7����oh�\\�����=̾T#��u"&��ѡ�\Ln7�CS�p!8�AD�.�nBL��&B"A6����
l�Hh��Q�	%r���0�	�F�$Q���q��A�!��#(' M�d�nH\�3n)��a�a�^HD��LHOFq�� Ta�$QF���.2�(�`�ұwϦ�2��%T%�뷨a9]g����'qOc\�+=����ۖ���fucU���/�p�9d��gs�����&W)�wݫ�1T۪ܝ5��CtQ�YV����]���n�1R1�aTf�HF��z��)� .���H��*Μ��^�*�ˊ\ɴ[�V��TC;��L��P���H�b�[��UR/ӄF�t9V廋/��Y!Qle�{�	aB�&x�wO��}�R�̉���'
�>6X~�?�C>�#��9��)J���fG�L�d`�x�V������=P�޻�4ps�0�vX�XĈ��4�(�$�סZ]x>_*�ѫ��W�U\<=�>&*�"%X�gd�(Y��Eb�@Q�U��0���6����#~�.��"�t�8i���^ď�XiTv�B˴=�ޜօ�ڒ�
3�S-26��Qe}	12�FbnMF�F��Z��y[��ʝ��fҺd�6S�#�N��M]��xP2��Ӧn�meX��+�u�k�F�e�A�RKV��C�����m��h�*iw���;���!B����~GʙtS!Bo��֛�A�WX�\�5�UekD�(�����Lj�H��si�*��df�7Һ��*�[�Ɇ({�<}��aR� ��{7�t�\r�cBwU��R�${���\wl,Uו�2��dB�Q��P6`j�	2T
A�"�v��ۇ�I��qi�C�$^�DY ZB%椙�	�����:������$�Ow٦A^L��D��rh{�/�UR��z���:������Ǌ�6h��÷�ە"�}�{��Xخ���0�oA�Hm������9`Q�ܻ7�R�V{1�`,�����-�)��L��z6v%1�]��X0h���$�ciw��7t�`%���^� �a&��V\c�1ٙ܎UlqXՓ|�WVU��,�=����E��şk��l��V�16�H-߫I���M�`�o�)�7���!ے���s��|��wΨ�ϖs��U��[A9�՟y�XP <}��y\ł@$|�A܋>t��V
n�����w�a��,P��VH��]�9� 3y�{��o���3�A՜-)gC�"���$��f9+���IE*d@�!�0��pj\���kP!�:�j���*���jܶ6,���Ž�����)K7�x�H�.�K�R��/T̔B��<3G��k���j9�,[*g|��S���He'!AMj��ݷ>��}�SSkf���6�4�ckuJ"�g�h'm�չ��e6���[���_%�u!�w,�3��� �F{�: �+�e�{��$���2o+5������<o}��/�;���U0�dCC�[�s�3lϒ�c�e�Z��+�	W���_eeJ����:؂Z�p�{j�q�Bh��,��6�*7��R����=�/!����b��=C�{D�B֨�S�*���
N��N��cLq�5N��$���y�;^�	b���8g}�μ�<�k�}�hԔ�HrQ�]�p�Z�CԾϓ��˩ʃ�校6E�#V�����ޜ�q����=)ӏ�E��Ͻ��fg�}���������
ܖ��j����������B�Z��Zn��k)*�ٖ~���f�|�׻������q�f�v"��H,&�@�Ŕ����U+%��Օe�@Eu���Iٌ����a�L|I}�˺k��0��}������of)מ��������l�G����T����𾺠�c*��"m�e����w��|4t{���cwv�Ĝ�Ca�--N�r5�{���a�V(	�Iy�S��u���э�,|�>�|�G����y��W0�Ʀ��}�8?�#	�B���D߶������3�Gȇ�I5!j6�	��I[�Yy ���362M�%;���-s���\Umkx�N(�����%�	��&c�N91�Q�t!P���(�Q�$�cϻv��)<�o�����䭐�"JL����n��;�v�0�n�mi�)�9z�m��U�����3������7X�3hU2IM����ڥ��T-�6�h
i����!�٥��]xE����w�*�wY��֪���Cjӣ㋷��:�W���L����v)B��1�\�𮐛�ߠ�#T�b�Տ���<�}-G�{��0,�ܠz:Rq�-��$�f�έT���K�z{ǡ4X��GbZE�tԁu�L����v��G˴9�}J�>$�(�}�+w�3��������S�n^��H�S�X2�=P�#a���J��F�!���=�g����1�6���C+3<�u����~��#��:���Gނ�J���6ĳ"Y4Ď6�R�~7w/*�R[��);�p9�sz�in���۷�+�R��$��P�cP��q�p�č��NS5���Pw��\s-XY��x
��6W@�E(�	�"�#�L�y��:ٞ�ϯ�*ƍ�W޽2R	.���<�=����е��.Ǯ*�0�6�/���~/��� ��鼛j��44a���ć/�b_�=��=>/�ڻe�C��y���w@��H�����@{�/�Еy]8���u�nm���T��ћ���a�S�q�-�����Tn�z��kre������0�X��#~ W�,'s~��㼹�Tp(�w��-��x䷝;V_:�W�9�u��YwNrI�;��:=���eCW�1�p${�>�e�Aπ����2���=�˧ʤ�p���t% 7%O^�~#�� F� l�%"Q��S�����ͧ���C�^y~Mv�Ur��N�J�1�H	bR�
���}��"����%�j��+��qU��-�5U� eP�C���!գZ����C�gq�gZ�.]C9��c�;�{���k�"b'Y�>����Pv$�e�	�UV^I���h��V�kUR�Ϧ�mƙLP��G0���#��IH%o�Xl����������=��s�q;b��	@���n��y6�&�$�)�P�y�'��i��mP�&���wkN-�9����rh#R@�h&��*iM�}��3�i�X`�������'�d�DkQ����+kUЎ1�"�}��͉��}����ZG�>�|� {=_r��oɏ���xj2E6���X���c��?wO�0�&�x�R�F��R�5!��~��&{﷬}�ӟ^fk�C��V�Vp���Țə�]W�ם�S�U��ԴCM��|�g�x�AB��ȁ��`"��B��{sl�Y��	Xef	xLa��+C�Ӎ���r�3��^�L#2e���ƣr37dx9[O���\�W���@�����$ƕ��cɀo)�=$�e�}t��4�B�\-�p���s[E��f)N�9_4�fb�x���>�+w%��W�Ԟ��e�m��B��WwY�k/��3�����
�%��{�"�_}�]}r/�����0�n7j^��T��~����z��U�e�V�1�O)I.3�����|��
����8�\h�+ү7�����ױ!��� ~�c����K.�}���	JI#A$D�
Q \�1M�l�_f$�A }�U���+\�`�}o��-�ؚmP��B��$�Q��D��0b%BBh�W��-�`��U��+��Sk�媔�gS�(�+QI��a~ � �z�&�lZݰ��!��Kw!������_ysaIww��[�s/�.H�6:�u�g�n�>��ɤmuk�_�<�T�,�����_Zu����r�"\#z�jD�-��O�]�_R�����`��ғL�l]�&��{�|�W��qā�if^��g�载���t�ۢ�#o�J@�������c��G��6Nc��x����ͪ��a��|=�xn������:�-�3)�kDSK����<��ٽ�D޲��!�Vosp��r��"Z�b��T+��V�3JMl���;9��[�f�wr�q��POpqn����P,�q�>ׯ'�`g����m�C�AE��$d�CaI_o}�3"�2	�{�S���x�p�*�1h�uI�((�)���28�O�TP�R2$&~�S�	t���
!�̯ ���DU0��D��8z$�`�ʠ��`v�}�S��u��}��6���>�+,�x����vc)`��;�� {+&v�o�V3:Ӻi�q^��3}U���+�����ʭ�!�媯��Cj��
Sw8T#��_]?���viy=��$�����x���ǽ��X�h��tV,�X�z_���?�P�wD�/^kUR�yK)����dw��2h�$.FCE$E3�צիV�6�7ޕMmL[[}U�R�|@�i)�uJ�HV�"ԁ�!�9��6b����¼0}��U�z��⃳�o��;1����G��s�!�����72��8�4�ܪKj�\�%�i��Ci�:#�n�V��)3etկ�]s�v��k��n����p <�+��I�ʠ_e��6uOu`.jX���t�U�7�@3^����m�r��	���l{��9�絀v�F�$�K�D!dE�o���isD{�*\�J�K%P�&����^};eG־6��Ri�M��g�n���;�p�{�<RIh���[lv)B�!����1ŜN��=�q*6�vQ��TnLP��̢�ܬ��R�bG�t����~_X���D)��dэa���r��{���g�E(�GZ�՞���<�}�{#=�9����:�æj�Y�օ��V>�{�UЪ{dl�]��.�]��d�L����i��&}ˡ�et�:a��ܬ�`���.ط����)|�L�B��>�ʝd�Ab>�4&��M��Ã���/t��hS������9��ٖ�9=����G��
�������u�5��g��R�w'q���w9N�O�˞`����b�k���Ll#H9 ��1�������4Q�ֿN���V{I�������N0��nL�ehdmr�/�fM���}�zU�)� � 'ވ�b}l�����}�o��ݜ{��%���ˁ՜����y�Ψ������z�@l��ߟ�U���<	�:���eW�1-Ԓ��ۦ�.�gm�]�U��_y�Y�jq��ĉ�Y�5��5\;jd���uI4f6�
"��/��*�}��mz������a#a,#�F#ʋ���uh g��]�]s��:�m��;��@�{?$8�{���|.��[�]·�z�p�Po���
4ga����x���A^�U�5�)�[�V,��=�,���S$��B�Ko����+s׊��AePf����T�M��f�ss�7��x�pҭ���AU��ʁ7	5$(�1���QD�q��E���(��rB�fHڊ6#j7I7QD�f"E�&�
E��`2���e���2"Ò(!bE)?DS`��u���$�L����D�@fd����S���݁� ����3��fe��@ ����$'���=�:�  �rHs�	�I �� x{���9"I"�I
bc�w^��D���ϭ�a7������*R�]����/����[v�^i}�ll��L���N.��,}�0=��PX����Za�vϺ=�̮�����0C1��5�b�>�	����SXRY�p���b֘��yɍ��l��ꪶ�D�*EQEE��ZI5$��!9@�	/̢�	FٌO6�)B�1[)�I`m��f(c�
�F�p�$M�bnD�O�H�i4����l�E���e����$e��**#J&2	eFDD8#.@�I"p�bN�p�00܄�8H���M�a �[$��1 �2�nAP��j#E�P��2E!��*("��e���tQs/�m�>����k��\j�����۝�򝻋���[�J�P1�7��n�6س#ޮ�j�3�Vv�u�(g�ZhiJu2�Hr��S*��ru�Ӎ�wUмͦwchaDD���{;c����طGc�.��;0���K�Q���X3q��!A��}�Q�ܓ�Ñ��8u+uY#Of�����V3V.<*��/uc*D��ѭ�k�>�[��BCcݩ��0��8�LYt�GBQs]tjy��&��n*F�A.%1HHeUA8�P�B�)��k��P�r�
��A>
2�H}

������3~�ND'D�T�j�] ��MROi�W�79@h٫�;��cf��Je!;D�Y�)S�m=��I"ݸSƒne	��a� !�! �:�ɸVbtE)n���������:��X�;�,𻬵x}bP`Ai���6�62*퉠x@�Xrfv��-��Hx��L����ix?
*R�*�^�,��|	6�R�]η5��/ևh�j�  ���d	�;^5AA������&��؟��Y�&ő.�hB�@|�\@�h+��d��O�Ed=n�Az�4���t�l�n6^���G����m�A�2_����@���"D�5Ùu��n��F�ٻ��өyi�h��G���
�՗�Ύ�ʽoAó�V�G��G.�D�R,�&�+o�Û,���a�;�����<�#���{=ɹ�V�n}�H}��T���#�yQ����|��(��q�ԛ�ːR�yw��{��3�ѩ5��ְ|�q�H{��_�����p@c�a$�D������u����G'�Y�܎�;���r��q�b�MI}��),�3zh?$ŁK$媤.c�>G�G�u�No9{jԯrjC��Op�Ǔ�0�)C5��Y�A�ѮT*��4�!4i�H�������P|�9%*�{!�ru����~�y�,��˸T2|�s��_+�����J���2@�5��{�9�y��5���t	No9�m�� Dng�1	9J
>�z'w{]�=� O��<�����j_9���	�z��0�/.|��a�5�'��>C�>���ϛ�����������}��L����(��'#�~����7)���&y����2�{9��
{��>�}���X���A������B|�����W�O����ݠa}�������ۓ�>�2��Ծ��k�3�}�RP��^��u�1/�����˸$)����gL�4�voh 9G��t�� �� <|$�L'��lu�wI���T!F䅴g�j�i��} �����ݨimR뻻��i�T��wDFx�wXR��	H\r6C�F�(('���Y^-���H�f�5�P�xK�Ղ��s������������U���#�}t�D��u]��^�s7a��΃p>Fs �Gp�unC�&����~�`e���#~4�,�QR�r�jNB�5��5's�A�r����FG��:�}޸������O�d"l;]2�py��@f׽�`6Gpw4n�3�%�G#�$;�G���s�5p:���������t�A)]o�~�w<Ǹȑ|����(7?.�ti�@y"d>f*Q��瑩�s�=-}z�/��r�/ ~�a�^F}g����5\��73�_`�~[�;�B}xT�M��ʐ| Dy}*=�I���B�O�g���.�;���7/]��q�b�5���:�����Ϯ��=���A�0���we��ԇ]`���=�y��B�{ֽ6k�s\�� :�J3�|��z���{����@5(;���
��:�SDj@����d>B��rN�~�S���:�]G�|������k���<�'9��%�3�<������A˭�gCR� �(Dr�|�{��9j@(�UϤ�����ݜ��5e,wD'$3;x}�xi�P��0������0ԩ˞��0Լ��������M��=�{H}e�r�Y۽�U/���!�}ʿf]�.Hxe"�d���ϑ-�`���ͽ�=�L<�� Q:���Zsn,rݺ��oD����
3�BCf�BR�/0���s��ps|d�T)�C�؇��yX=������y�!�dezg_3~E��9F�>G#����a��縇��pw�!F���5 �9�'��.��5���$b>��I��{���5� �ݳ�(�Ip!xa}���Dy� ] ���/#z����y�5a��=�PП.��X��0���=��|��!@����de�0��:����� �Bzs�=�@��lw����AA�h䜺�܇$�>I��49{�n�;�2�y��s��@u�S^`n_cr?'�a�����3���i����ߚ�,�ut���ր�4�����#�P!��]t/,��2z��{�G��xgXj��4@jAș@CZ@c��tUfOup]�@���� �z�������vT�.��������N����B�0���fb�"�,������?y������fA�wd�S�y�1>F�E$<(�>��>�zm�TFĒI�V yU]�}�W�ZBnC�qϘn^����q�2�{��@�imB1
#�>�5׮�݁��9�ߘ���<�y��@e��C�3�$d�#�b�x�8����Kr�;=-� 7�5~�b�U��=^�ox�O�;���l]�&��R�yL����y�}S;�wV�1�=��=RQ���aͅ�V�}�B|��5[�=��w�d���Ns`�QH���#��-��P����Ȣ$��Q�L��vmK��I�\��{�Y P{
&��|�1�CH� �S�y��~��ԗ�j��Ѹ�'V\�>N���4z^{ָ|��ά؝n�pd}
�Nf`���g��z�oS����Fb�j� )�i
R9(��8��fy�
����UO��"�u�j��)���1��b��Ե!�ڵ�$�!�05�!��̡�fK�ԈH_\a��	�rn2�[qH� 3��{l΍&�EZM��h�����?Z��:�T����,�/E:��s�/�����axa��ƴ���1b�0�}��b̗W�G�K�pI#�_z< ���iUO�,
 5<� O�?0V�8h����M�otX�������f|<Hm�U��\ (�0�Z 7sX�o�4d�Q���v-�Y�w���T>���E/9[e0i�5�&i�}�g�Ft�[B���3��S���d����(v���m�yJ�l�����3��J�}~��qS���!]֎|=�?���Z�dw<�%N����p!�����2�(�ˡdp U�� !�2��;�B�ʘ^#����L�xʎ��j��D��pJ{�#J�H,G��g��.�L?��-�9�;�7�+.Ħ!;���1Q�!Z�|2�N�T
��	emD��w�T��k^u��z����Wo�>t&���A�&��f	��.���)���g���ҲU��A�X��oE��<�HB����;��=� �����I��}���l�mq�?]\<{���|�#��Ϙ?U;�l噁.��0�:����t;���`���#����q�$ A S�=(���h�KAA�i�[� ]����<<�j!)�e��A��Q��籱�����y��QGԐ�=,h��4�`�~ҿl�%�|�[e�bR4��m�@�	C �����qɜ�a$��$���wRn��6ѥ,�˽��Q1Ɣ�?1".HG6��u �FH�Q&̅ dN):Uw;���9h���8`T����-��i�7���3��
���Q�=�ul�q���2	*��Ĥ������29��z3
�,K;Z���q��6�cC2K�g@���;AYX��\*�����W�C���:���!?G�*���*� D��կ�`X�F;�-6sulG��:- E!�H��B+2Tȃ熧-��t��N�&�����#X�XBJ�@�Bt�*�,���ٺ�xf'�f�D!��K��X��e�`ۑ�,����oGouǽ����C(R�٧mZ���!��\��񙁣0x��6�A6SK!�#`S!:Y�FN7%�\x#Y��W&n7d+y�fvR �DFV�[ ��ϩ-�X��f^S0D�Н�y���7C;�@���EW$Yumq�44esfݪ�@��&k�|����!����:Wu������@S���d"�@�
�ٲw�2�Ҙ�.��u^�u&����i�ogs2u�N�R2�
mC i@���# �aK��H
��U}م˖�&K��}��9A""!&e��u��m,D)�����f��ӌ�g_!ZBVN������uxxe��E:J#a�ɱ��dsl�+�wB+���$�F���c�"Ј�R�(��<;
!�`YkCm�OFn�����4pO/:�hQ�U,�nELp����}F/hʁ�b+X�xDl��H4��Y\f���665ω�5Y1^�f�#����yn 8^��F�Ì!��a�K�EC).D/pٜ�����xg��&��c�<���4o&��#5|���!���iE���4���L�������>#�@��* ���oQ�ȸ%5���.���9٭�@�i%-����3!��K�i�0���6�j�!R�C��[�|�{�4��Gf5T
��	e;Z&r��jʂ�b"[���H^=mP���ؐ��=��
P�$Y��3δk��epkb�bך��5��H�	=�c*�����;��ȦC|Wg.����k���+b-�i��#O`��D��$2Li�՝<=�~⪟�����4'0����Z�]��\���xd�z[d>D���H^s�H�#2Ӽ�7!k�d>l{�o��<x��R��U#Y|�͚!���/,��]V���<=ᇄ�o	��V���$�.DfY/�=�˾�"��󿯟Y�9��0��$9 T\#��m���PI���i];���"S���x������+��2$�M�5������ ��[!�B��T`\ޮ��iϣŢ�a,����O���a��̰R��%��Տ���t�1��@لIZ��� a�N��S!E��{��[=� ��\�U�dI�T>����⳥�.���+�x�h���{�A���uԂ��.�Ѕ��"���ή���� ��<�z�����s�ۻEa�q5E�����̉���|H��nk��`;? SߟWc��/���s���'�u�>����퍙�/�~{O;,��U����O�[�]♇o���69=�qOy�}�!>������������/��P��c����O{#mЁ�,S���U��X#���������ƴ�A�����m| 잧{m�{��o���5���	mu@���;�9Nd�|<<� ��M��$��F�(�߯������б���@��7�y���s�����zm���"����9*��� bE~���ź-�e��IPs�'�(�]���Gx]�ņ�eԧ�rT�mk���l��)�p��9��q =�u�SH������R �)Ì��8m2�٢��^庰��).�Ͷ�C���f1�Q]�/��Z|<2�K���.����$Hmp����l�s2�Cz+V��_S7\F�0��)�3�Vi��ǩ"�[3Ϫ�u]�:���(�4�vX����GPD�Й E��5����/Z$�i&�.2�n(�9���4ʎ�l�<����	�TK�O��������R�j�m��Bd,�F��&�M�|㍘���4�!�L�8a�eL�y����y t-����q�8�Oz�&wU�[K4[5$���ٽ~������v��c�%�"E�4	�C���!8T�\�E����,�I!�7���~����S����#���S"UY��>��H�0�l���Ӗ���Ef�q5E�������b0���[&n���?�C��43GwմJ����*$;s��8�����	�,|=���T�f-�G��@N�d�dL�U@���\�;�ｃ��>��o�|�"a�A񃱵8�A8SC!��`}圶��h������EQ͏11���-���j�Hp]�ͨ柽����aDD�7�E�-�e��IQ�2j�|�������?T���X��f�j�`�1�(K �n�u�դ>���+M���Xr��vLV��o$�Z�C5�UH@�E��FG2.�� ߯��4ֆ��A�,<<^*zh����f�V:c3�yGN��>��:..t,7'���Y�ћ��مڐ֕����%��H��`�kUOUX_5��42,;���j��9&h���%誒�H���g}k�;�3�}&9�z]��50�$�����f.�����kߝ����n|�1��虄����`DT�b��s�/s�f|����9ST�D�M53@$����_�u�f}����+=!Z0'�_�=LSy�k���5��Įo}�����/�>��eͬ[��؝���!����pXi�O���~��c~ܾ�3���B�O�^T���C� Ì#��߲��7�^0���Y�
qc���`��ˮ`�=�ݘI�]Zz�!�W�a�� Φ�(�Jj>H�x�1ؽ}�H �Y��klP�@�9S�y۝Y>�IV��'O��0ּ���||���F�}Gz<N��:B*���޽�4I����o��P�N��)�M��A���y�o����-B�=�:���opl�91�uGWDS�dQ�/r�UHj��r5>���z�ЏXf҇m|@��|�L>kL�H�D��"6���de��v}�t����͘_0vԂ�;�������XJ�{���?3͡�k��Jݘ�.�sHJ^��\LN��dw),�J"���õ��2���ؖTx�߼/�������|�\}�8���w��Ϫ�Q&�,H��%����	�2}�����S{�$�6܊B�ppQ��݀�ݨ 3$n��9�t	ʷջ�]�ؒH�� ���Iy_Wn�UU �H�ۦfqN �l��v��S�ʛWQw��g��d����J��`���]n>���;�==p�]x�c�\��rs���H$b
�<�Yv&f	��q������e���j�G<f���9�����B����pw璔/�D##4�@��s��̱��u�]i�*/e���o+��$��2Dr��kn��_p���t�Hj"�o���zP�u*4S0�ۍ��M�$1C-Fdi�Id�"��a6F ��Mȑ�9�dd[.�Q�� ��$15"��$Jd�7��#(��4�"	� �%���-��p"LF`e�܁(I�B6䐔Zl�J"�q�T�:�h>�PI�ҡ�{��RR�gT;;lv;o��}�/���sa�u��*��eS��u�����rŝb�;��]#��N��(����=�JԐMs&Pn����>
�1�V�o( ���t�Ln�U�:�i�ԫ�b�)�y�wA��S��+ti��m���%W����ϋ�~E�� �h{��c@�@�ߟwb�o��K�CȠ_*�a\�F�W=v)l�s}���� zeAdV�J�R��xNNŊ�]3KX��T������콋�P�M�c��(V�t���#AiwH6��<O%�G��j��<n�-4����1G�V*���b��r�m�!�7<���JD��Se�M��? *�5
m�����X��,��6'��kt`[V�]HW^B��(��R=*�� ,��@/�a6�j���y�V���Q9uN
�����a4�Ψ:)a�=�xi�KU���}3Ek\29wA���0]#9Ң�F�p&F��d�T}X�M[�N��iQ�`q��$�H@��� e�QT�{�/P�df��N��ߗ68�z�ް砀�A��|7I�_�EJN��ۏ2���X���.�[y��cZ�c�/�*��Yf�5RA*5L�!4�	���F$2���];2����ۂ�Z����q��@$��$��u\���922�w�YCߧ�2,#,߀�k3�!A��b�rX��<;
!�O �����<����ś(Pnp���rɪ�R��T���`~
͛[�� �~(��FT�d*��d�\++%S�������ޯ>jTע�����K#P̂NW�"m�+_��~�̻G�(�
����!{�_�L
e��ƈ�x��ʪ{٥�B��0}v����g)F)��'� +C�m�}�������'+#�%5����ӱq!G8ɀ�I��L�L�6p[�ή27)2u�!2g�;�_/�W�"|mh�ǙC&�]���-��Vyz���NJ_PM	���C��z�� �M,�o�`S!:X|h�SԹ{��\4��ک0�oe�C�IR��/I��[ ¼���k-y�{�F���͹OW'�G�XӜ*����s�	�dD��¾� ������9b�I,�.��I�t���ٖ�w˥V�Kw9���|����K��V
���L$�=��D>wW�۽�g�>�f��o�tW��@�FǼU#���^�M��<�^U ��CWs٣Z�Ak�G�W��?w�z!Ȱt���Q'� A"�p�##Y�z�'"!�Z��S8�1�;1�y�>��S�5�;,b�t�E�`[/������w�V?v�:X&�[2O��5pI+�J��]��e8�M���z�����ǒ��{��W,�[[a�!�#�O`�+)��ųM]�2>���O	��ND3��@��w��p��-�������V��0����{"��L���L��S%9wAȬ:�>���>�����\fa�!8ƥR.���zc�3r!h��s�����0���\�i���&`&�bʿ�\�����]�"ר�>��M�P|]�ѿb����x�����͔Ĭw8��\��3�ojL�7o������z���&+��7�7���ll����H��Ub D<���ϯ}����_FFC����m�<�;�k��4-�(�?�ow59π��unS�hoYf���H�a
0� 3o�����T�eԘ}P�m���y�t�qP)��n7��Ӻ+�&��`��Lm�~��yh�ը�k���Qd�a��]A��[92$�*z-�tGt8�SlSӓ`
�\\v��@�A��ĭ�k(ړ�Ѕ�nF��7̷@�<� A>�a�Uִn�O�E�Hivj�'1\��ٛ����@ �JRTaR�)�xvC�F��Vv݄��̭�ީ������Z�]���6M�݆�4��I�4�бLQ�bT�����;|*��b�_`Ku�J1S�EXY�ć؉l(;�R_�F=����B�/Jr��J�s�b8�5��^����VM? �6 �[�T�����)Wݖ��j�j�ZFC��I`!��1H����l��M��p��U]v�Tq�Bb��Ԏ)�˖wM0�.)��"HEj4�����n��[~"Q�D�,����'W̵c;T��u�&���>�,W�FǀPw��C1�m]����{���-mR���n쩑�N[�*�9����gD� j�r�f�oH���b������+��'A� *Be�Q{��l@�5fd,�FZ(�'84G��[�O�t�}b��A��QYM���x���{��U��D�3f��a~�D�r�J��돚��D�w�7���= nY���Z��8)��,�9�c	\�u��ƻ;��
���ܜI����3�S22!	
">��̋t0[4�)��3s��#	E$�(�7�"��b�n� ޣsY�qc�3'���w�Pʷqx���6��v�P�}�R#�Q��T
� �"���d\��^"P�n"N]�H!�o�����H��
���dr-N1�/���e���&����i�cd��3�5ٙӟ�&}ޟ"πC��c�*yY��]�v���k���(����pȃ�n���~�İ�E0\��D�_j�d�H�Ϻ�id�UmT�p�Pb"eL�ə�q'c���]n ef����,���><1�dRP�)��D��vI��gIp9P���u��$�ZTQ�~�jE2N��Cf춌 W��.���Vf���Ս�$>�Ud��AL�"��m��G��e~�q�K�I(R�B����G�z��veHw�N� 1��4��򪃑W��MQvtM(�0�#�Wh�Ѿ���Z`��r�M�E�)�e<������KZ5^ό�%7!3a���*�D"?N���۷��s���&����[]���.�Q����v+����wܝ�Ô���)0NS�|Cy�C���\��%G~�11��KVІ���#ܧ����i*����A�HJ@lM�١n��f�I6�0�J�
�*V�xx@����φnCO�י�hV!��{4-BvT���݆�zq!�>ļ=�!�[ؖ� .�F��*���~'�d���̗o0a����ץecFZ�ұƻ3*m:p��Cҕ���p��B"{����9h��9������--|��Ki'B��` A"H��##���VG]^�V �:���2�A��gD��/�/l䈢�x?R{w�}(6S��H�Vk]��-�tS]TEM4J��f_{x������\bPQFnѕ�
jy��]������x7���>�Xvć犬�@�h'��S<d����UKv&�`y �
E@�jn~ �U��1J���/k܁P)���ɐ>h�(*|�ڷ�9���tB3���1�N.�t���/��:�j���;� 1�B��Q}[D�����F[)��n�'�x��q�~���Fӄ��`<�("�l	dNSU@�����8dZ*"hȖ.!��:=9BA
�`-��dKP��{�[k'Nk�	�P0 �R�����aip��$�n
Ԍ|�ܷ\�~�}���%�A��3W*AF���	�w�g�nme�r%Ky8��U�IihS�q
�T+�dӼ�������� ���c7�bg11�OvF�ѧ��C���/�� ��V�]Q�d[��٢RM����C F�����Fu/ʰS�J���j*��CW.�����E���Ǐ�����D��������uD����`<�'�t8���Fb�l�<�R�ٜѤk`���T�<<��.�ﭸ�9�� �!�i�1E2|�.,vNe��L��Dc�~�>̫6����$�~��}T�u�x|:�J#���2�S!MN�(����Pr����Uot� �$��hH{x��H$R	����1�E�޶�t��{8�����a��j2W��DE�YV��O�χ��!}*\e�vtM.�0�!8�tT��{l��\��v�*����8��C�k�.�y�nH"���14w`K��S"\m8Y��"�̶ћQu�nwUWU,����)"����% �%n��jm�M�e��(`P�����L5�\�ƔKy�3z�]j.��� �G���v�
aQ6n�-g��@ C"!�f����>8���5�W��]J�� ������/��C��	�9�S��恶wIِfv{��@V��4Q5�$��W�M?D@��˽S��^���[�S���z��G�xS��� �D0���9�)���f�]��� @z�E؁�ʹ�cT�a����f��bg�%�	
0@ڏ���{��\���Y�P	5� JPl�2�#�ˁ;>����=�}�7Ӽ~�;�NvH�o�x<�?��c�(k) �x|<ݒ͙�����z "J:���}s�>k�y�ˉc�y�J�Y�;�]����Ǹ �	nc ��6@�b�	��C������_xT��¹�}�8�d�� >���*��S��z�Zz@��OJ��{���AA�ߙ�y��}������uOk��Iv�;:"�րȼ�.}�H�/�Lfj>����5�A�&��޷;�$�P�tDH0"���&{�E��G��k�ێ�J]{�����dPhH��u�U����jwU��R�${����z@v���	UA/&"*A����p�
2"ԑ8Ph�_���C$T�K�����`֖HT��l�$�Qb��Ӿ�9IC�^�~�����^^��'��]�p������rxV���@Ĕ >�K��[
7�ו#�Q�L��d@ce�i����T�=/�w��.�������gD
%0�4@� : *^��@_E�{�!�F=��x�\
��$wx:� ~���𻁲�q�@\U�������d�1��,�q�W�M=v]�.���ᒻB{� =f=3�|6@Q,�>l�k��-�W;F2��z��k�A� ?�� � h66['H� ?�K��e{���^��~�k�1��M��P�����c|�I���@^�8�gg�������Tא�[Đ*�2ޏ{��D�e����Z��/��iF�N��9����`�HH�(8���4e��Q�݃���I��(w�ghw&e��JW�j�?��x�}�D�C���o�O{�@<@)M�M�*�%t��a��'��ƹg	�N�����N�v9�y�s�6��ku�tr�B��vaݺ�9���f�^d=���ʮ�����"���+
h*�U��ef��OT��3����{��ز�O<�6kb����#i]�c�6��=�{��q�21��m~tm-3N���a˒_��!X����ܱe����&�?9]A'�V����T��)ygx�����8�S/E�ճ 'Tm�n��r�AW�8��.���r��VT6�&�l(����¾_�,�<o��b*Ъ��������K��B�����h;�;?�����G���'�]��|�^J�������f�x >�=��
�U�N�++�̳�I��A}S�� |��qg�l��{�*e�_6FȦB��֔]��͔���sP|����3�<R�R!!)z�m�h�n�f�I3�|6J�s!�H֗n������ܠ��;;��!RN�#AS�����',;ޤ]:a��3u����oj_�Ӓ���N�:�NP���7����N�\��������rs�E��;��z�0�>�讣�9{'~e''$��I��b�^F�� ޺���ZP���|`֮��lyD'�@�&M#��U�TóV�c�b�6z����҈i�CA�{�9<W��7��qC�|h�}��˦|���ro�/t��̎��2�۬[��2�?z
���������B4
���T4)����;۫X�m3:����F�8C�w�&�䬵����>@6��� �:�A�k���>����׾mw>ABn)[κ3�L��y�}�(|�Kw����[�}�����<����C��ef)����ʘ�͡j��<(*���P$p�ޜ
�m9�~��u���E��7�Z��u`�,�c㳛vR�����"xh��!u�����]����[1f���7�!m��t5Yf^Uyw�1��E�6�O���FGB(؉���!e���(�Q�J(�a�-��Q�c�!J(��G	.9n6�I�CA@��0��F7�2�%8���m��*	&X��<�߾��{$�L���wv3&ff�|8(��{�� v�v{���z�H =� $�'�������]���������OI I ��<'�'I�I%�&|h�^3�'�he.`Wj�Ko
:�4���Σ����n���O;B�Uz,������U��$��H���󱒍\��q�@ugXD��JR�>C�Y��pؤz�|oS���R+�����-���꿏{w����k����\�(��%
D����¤���0��i8��l��h�bI�H-�$A�Xi�R��ҁ��b2X��Ą�M"�j`m�2 [bH���Q��I������IEfz2��1I
�1���L��)H-��i�p��NEiƊm��l%(��N'#$�څ��"0�B����)�#JCe0�����"&(�d���'��Q�l�ͻ�`�tF`
fnp�PҝK��R`�c�bu�q������G��=#�Ma��M��v�9)SG�Ճ�9���J.�ӻAGEE�U᎞M�5T���L{c�D���xҌ
cof�/Ah�W�0�2�ʒpշҌ�\�G����xod&�:��䧚q]gm�~��TȸI&c���+Y�)��gVW� �:����FM
1iՊ3�fi�RRyp  �Ѭ�0��g�4�)��G��F��>xBX �X�I���+�s�+V�G�1_�9mDM�&���	3�ac�0qQ��@�e����G&���$	$��G�/q豘��Y�zmG(�׽��ZY��۔��x1`�B��eJ6�[��n)��ń�q���k�@�	d�`�y/i�B�=G����]��V�Y�gp�n՟,�����/N���pe�u��a��X[0
�۰a(";:��)�O�gކ��O`�B���{'E}i�;k�-����ckc��ԣ]nԜ�A���@��wG&2¾���E�z�%���$�Ǵ��haxaٯ����Ж��/
�^�S��y)�5� �\��Ć�������,-,�A
��f2!�>�{�l�Px:r0��E	ɹ�%рr�\�5���m��|�p�m�ՔmN��B�Xw 4��z�sS�P�A�Qsl�Ʒ@�,/ ��3�MT��b���U,�����L�\�{:�XYMT�e�_Pִ�	�[]j'u�*��z�����`���8��o!�ra�NŞ	J
"N�2�S!MN��툯��k�x��:Q��tm(7N��\��$Z	��\3��CVA�o{� F<����]H§B����=�]��;�o��> yم^d��^��S���=!���&�q���1�������;�?��g��*�x����Hd
�U�a��g��a����� ^�O��[	�	���J�Z���

Q*����!� D.4�����i�ߖ P]Cy������#�
?$3�h����q�ȁ�A��T1;�#c���䕵UB����ft\�����^�����|	%� ��!0�R8A��#,�č"�HLM� I	�5�fn���K �^̙ܽ��vA�Z.�g�W%�� �ޣ#v| ���B��b���}�߻�\V�ݡ0�bI$:��3���:�e\��=�`�	��ަ������惥�-�}CZ>lR�Ɍ����Y��;]�c.����r�$�hFI�{���98C`�Q_�h�h���ؙPs�<Gr�G��=n^�ӹT����5Յ<�8�D�U���|X���Q�t��`����i(O��q������O4��5v(Vm�4����i`��=f0�����Q��`��Yc_A�i����k�f}7�3VCT�1�=cz'[~q�\6�i�Ò��W�eH�Bi��Qk����K�a�]�?�:�V�ؗ:�97P��L�4�>�>�e��B��0�,���~�j���N"k#��ON95��z��� �j5�W��\ߞ�uo3��s�u({�舂e�)�$�9S�W���F��>�\��,����]h�l-ab���aN�R��5W/۩l7��;�o����4�Ls�>ݱ�]Q.SKЖX������%�[&�a*;�U���bv�&�s)���z�%�3��`��4�iG#=��H��k�%S��� a�^6ʇ�OH_3���L�M(90��Xi��{���go��H©����z�	����t���K4�M�OE�Oy����~Ba�f;���|�dIBq��W���u�͒G�  ���������$B�S�
�ad3t{`}��f���cD;�3`���٪U���lڂ�!�#��v�6#�g���}ԧ����)�%��bD>���s64���P޼�I3����l#m���.n=���9�(+�gwt쓱	훤�G� |$�$DY+>�� If?Rym��)��C�C�d�d���~�I>#h=�������ȈSF+;f1�"�+�����<�<��1G��TO=+?��=���5n��]S*/�0���ذ�3�x_�����>6��@{ȁ�<��P!�w�{6ʹ)�6�D���% ��ch��%�p>K���	����qQ��)	�ꪀ�A'�BZxpي�f���A��X|22��DK4B;���J���]voOwe|���C�9��ut�,�"\c��6ح���꘻s�����ҭ����1�=���>N�'�k�C��k�+����B:�i2bԑ��1L�����co?��sՊ�Ĭ4�X֓��
�"%3��� RYWoD�䘰IlB5�9���� P�t�H�rz�>��37�ev}����u(�(����gv�HL�r]q����^V����#W 'C����>�d��?!T�n^����"�V_����־�D�0�*�xIcQ�����X�;�����C��r�	hP��hq$5K�n���"F�'�G���c�ǥ{�.�'^�=�**�FI��xY�B�ܳ&{��gP����ݒ]�I��w��
��Ojvά��D�JI��xx�\�`��@�.��(�ĒG�v���� �k�|��4H��r�Ua������m���AS-�F+9g%�1ʕ��.���`!.�*I���C1����D�n�\�,���3���		�i�DĂ����_����Z�T��|t�*.b��8�e�Dw��d+�e�dPp�?u�a���q�6�AdJ�+~g�	w���9��C0v~[rۜ���i�N�-���ZÀ���G�����L���"���2oS��Wy�< �� G�#�C�.��R�A�R5a��>4���=����� b9�L��Bv��Vc���]K���y���\����=�8�����b���a$H� �ù��}Cܣ1��y�Q��@��^�{t`Ux ��QFE�����md�'N8�J�`����./�L�ى'�H3��y��Z�M唂��Q�sc�4���fO5<�p�6��,8c�a��&2�fC�<�ʮ8V���F*�Y�BF4$X%� -��QF|�h0  ����o.5���e��7�LZj��DDF��Dp^i�%�����,�w)�LJ6���������QI,m2b�!�^�
�������Q[���E.�p��=9w~s9�8i�6�l�3���J���L�Y#��2������|��w�`/ ά���.�U)�z��wV�od�����=�BCvk�4v���}����^|z��g:������۱g�`�'���M��b�vgy�@z��k:�9-֢�:�� �o��m�!j}L��Hy��Ƃ�D�G�f;3u�eO0��d��-%���I���Jm=��1��+�졜�a.f	g�#�x���ʘ������(���u�M~�|�a�������u�E{ח����DSD�f'Pϳw2fK��I����;*-�'y��\k7)�P�t$$ƌ&9#�B$Y��f2�%����;�M{v�u��ZE��+�$�oK�4
�Vh@���)z�N{��4���T�e��:�|��+���M���H����W9���)���B���U�Y@�Ò�4�mN@���u81��X��	"8����'nU���0	�ި,����FQO	-n��ݝ*�`�$C�0�N�2�H.!*ض�����4\�
�n��ᤃ�*ξ4�#�=��eX���	qZ�I巨(EGPk���c"�]!\��꘳���e�I��3�U��},�j����qF�� ci[;�e7R(2���З2��� ��d*:A�{��@����!H�f�a�v�D����$Y�R`k��2�^�%X�dQ5��=�K�6j�m�x�A4G�]�_4v��O�z�=�F�Қ���%��-[��~���]eM��XO9V��wdc��M=���1�*Ê��j~T�{�U�+�R���h�	F���R%���P/��2B!�F�
)IDDi���;�[��k��e0�u>.�'�k�DZ�Si�����+�v�w���?2�B�����U�Vy,kI�{{���З!����I}�rq�B��|Y:�/2⦭ح���vM$��;3����S1=�_}�s�����L�.0w�����-�%�Ω�*�e�k���ޘ�7�ܯ^��jl�vP�R�Y}n�D
#,�����9*`��Aj2�M�'L\�^A�.;!��w��7�9��M�ATd�" %�K6�N3��T��I�ޏ�K�!ck� ���(�K���q-|��P�<]=�|�5��P �O�X��o�����	�A*�jk2�+�9�>{��\T�b��%��Φ�F'7���/��P�S#@��K���nT�t6=�Nq��XRYr:L8��rF'�����aÝ@Z�]���)g�s ���O��ze�]�?0��Hn�$�R�����={��\A�R`Ҹ8Zv M�dA������fb��8��)��>kn�Ƃ�R����̖F\�>O��[x[
�bZC�mfl2OD\�"ְx��M�$A�T�����v���$��.Л�ޫ�-��ĩ	���:c;x� ��vfS0�D�RC�a0�US��K�5����U�.��C�%�O��@&�B�6�k��m5�כ�@ �0�*���:���Tu\fj���c ���|Nf`1��|o}V���8�4ZxIsi�v�V�=кȪ�PH�l�� ��,̯S�'� ��+JU��M��7��_|6o
U.�2H#L���\e�Ii�O�W��֕�I�Є�&��9u��L��#V�.z��2�d��D��i!-��-��lCbD�i"Zl�	E��e��y��;;y<f����hj(�&r�ɻ�c��1f��P-��i��$�T��!@BDB���Z`���!�ߘ�֧���ձ9 *��9�6�G�܋P�Hk���ep�t�`�cG!�ɋ4$ǹ���n�D��%kvJ>i8̎�+�7-� ą�q=�����Z۔�aD>6�d_[�(���k��B��(`���cL�akYyz�
d�Cچ7r�ɪw�^	�΀<7 ��
�!��TB9<�Db��\����M�{��%ҧ��ɗ��4�E��N|ő/X���;���=��>����J6��͑�(��dx���+��/��䗼 26���hƩ"b�b�{���W4n�W�<��e�M�Ck!óɀ�ZR�s��������W~�ÖPm�T͠ǰ� bV��	�'j�U^;��9ppތ7���Q&a�*��*��%zM��̗�L/�t�.'�c^d��ըƾ,��[���Q��la�\4֪ީV�ʘo�֝k/î���*U��*K�J�����Y) �ڂ�Aq���Ι�=u�h�V�;h>��>�Enx�U����j|6.HʍM{�\3eAVP����Ӭ�R���E�얤 �YV��k@ �]6B��V��+��Ai��.:9�c.\�
.������A�9����!�kGǰ���ض����y��i����lS&o-M��L�L�K���a�=XY�}�}�����e;����2@9��k�4���ѳ�\����&�����";���P���N<���5�6��wVGn����v���X�J���0jv�w��C�׃)��Ӽ�S;xj�a�7Wq}���~a�RzA&B[�)$�J�"�2T�H��N#H�#p�$���D�BS��|U=$�'�y��US� >��ޒwv9� fd�zHk�@JZ�wcn��$�U:7wa.��n��32@�r����� 7wc�n��>�� �f��R9�UfL�U�q�:q�Fؕ����f�Z�7��wZ�A$��������g5�WϋF�e��z�T�n��OGf��B�݊x���aN{���ۓ�R��c+wT�е\{g��ح"���6��K-�$�0���|N����p_ah��:o��S�5�t]�<�*������;�t<�]��L>�����mEe���RB�0�$I	$��D�DF!RF����8$ ����
P��!m9!I��OH�2��p��*9��nBahH�-��J0[hQDp��2$сL�am8��h��1��%��h�#.�Z��������Ź{�����4p8"����Jp����|ˉ|;R^�D��^��2�!�qrgw��=Q�J��]���E�����mpFFق�Υ�5�9�`D7�(���_TG�ّ��Ӛy{��Z�9���{��9�n;�9
	��mYR$�PY8mf�Z.�ζ
	J�Y��s���|���Y�+�>��C"�#a8A]n,�R�G��6�!�%��
.Z�Uz�N���>Qi����^��s0g0@qeۧ�U��4��q͈��ZԨ�?L��CI��U��d&�n�I�Y" -��ͽ�)Z��SE:$�}�=���7�D�(<�]�����`��;uU5��O}U���Vu�S��$�!3�7(mW0<�Z��r���̪:<<a���}=0v��ǆ�&�76�b���t�Z\+tP�a�YU�z�[MmuP����2��]Z�Bj#�U,T�2��{H��F!�t���[X�MePkD(R�ՃfA�v������`J7�9i���U�׷�-�#�v`'6}v�]Ap��Ž	Y����X���>*���1�nc�F�ڲԃf��mU��5��rC�X�7���q�kv�旑�y&��.G$��SP/Q��WR�����rw�5.�F�{O�ԗX�"�w����`� �	Le��G9'eE��t�/+M��H�+��9�лdxdP��v��J�c%�^� �$1(e���c���W���a$h��ƣ&$���v{�r<=
�ބx
3��϶�E,y��CU����*�Ht�J�^X��sM<5�!u$ׯ���ke˸"bX@��.Ǉ���n.��{���������H\n��M�nt��vD����9,L�M��wT�Z���<�xFe�r�����96������˴Xbb�R;}8�3JL$��a�~�E@�2�>b˺"�
xSG�<���l$��a�h(�epU�ul@�hSL.�aD9�� L�}v�TE�0��e���]��H�C���1�4ː8{�g���}�|�8�	C�&ER a����L^����>����ꮪʪ�^8��K��3������r�YY]�u�>�gw��#=�:�{��r">�bG"TZ��:�@��z���%��1&�܃|�j�ֵ�	i3'*�fςu��� zrJ�2`ԡ��1L�����7�Z3F��oN����X(擒��"%3|i#�犼ޞ����%-�y��73 �ތ�ϰ�dDœ��&e�nx�Gtl� ��a$N���Mɋg�\���Yi�f�y��"�����0�����0��8$֡~JSM��NǚR�`ِC�0=���(Vlt��<׊�N�I�~q+]C!�G[e�g)""Xw!�0ue"�'_O؅�C�j�(�6n�Ȫ���2Nd�-��z!���5q��[9G��-����r������B�8�<���|$0g��&��x�#�hF�(S����΁��r���浯�y��o��"ACۤɧ��~{��{�b����b�o_i=B�1)ۅ�7fr�VVVrm�
VD�!'� H�E79���Xg0�#�Ѣ���*S�ȼ
E��V���ܥ�W����6U0��A��5�D��dp7:U-�{.��L"���/DnU�۪7���0�7a�|O� ���TE�`�e?����8L���YF��!E>��B�a�^R�B�R��ޫ�-��x
�|�֯T֔���K���O��s�XDD�c�$I��3���5=�����B���U뱝�e�A�$��9P8d��{�pl�t�q$H��<���3W4�Ȭ����e<D��H�(���.(��Z��=ֵ�oFAnD��`)���$P��]�7��R� ���\7����a��P��$D���$Du����-������]5��*7T\���.�jY|R��DRR0K-I
��J-�6�st&���+��I+IF%�;&�t+*Y7(��j$T(&cj&4�p��J)!"�PD,$�q��r3!�'�j����3]WlQ�N��r��(��@��˚��%�|@�QJ*S�%[������bw���ﵭ��(�6��Ja�gxzh͂�9;�Þ��,ND�5����kҐ��_�=��(.m.՚K���૕�T<q���1
�9��b�$����C�����x�9c!�~")Q�	+9�Z`\�
B"eQ�~�Wg��B#XES
i^��k�w�����������Q��+S�*"��<IM�VKI�ӑ��ڏ��E�#�5�U!|�����m�A�A>���y�jX���\4�$*ܜq0��*zY�pxx�K���Ee;L,1�9#�8TI�8�7O���*�����Ā=�^�EiA�@l1�)
�Z�6�֔�@on9aԯ��������xId~�$�x����Z���o�}��-I56
���vZ�V�s����N��s.TX;��l''s.m�B��#14�	&�&�AyȘJFZ�G	e&;w/�pdwq�;�MR6'�e6+���-$�O���mG�M�4�7v�Q�K�,�C&-�� �$aHmmE�O	-m2`�	��;�X�����@>e��W�,���*��ؖ�b�!-�y�h�op���ݜbTȇ�U����>�I���}w{SX<� �ZA�����1, [\b*堈�g�交(q��e��"#z��r��#���7K=s[�w���˾�9.�Za��j�Hp���>�<+_u`��� c(2a%��c�䪃B�bUBg�F�G[��qH�0
0L�����7�3�V"d���6�%��fd��L����EҶL��3�YY�z�$��*J�#��v�������55����+	�Q�'%N=b��y;uK{\'���������}
���Zź��QS2�<����w}w�H]�j�n��]}��vg[�]a�c�l�1��	�2$6 g/E?�����1�� �9+,���">M��;"�%��c!��}��6i"�z�1!�4����e@'�J�m�����Ob���bԛ�F�6��O2dA��7#�=ң�K�#l�����8dϭ���s<k~��B�����u*�cY�(���e��C�*q�Kw8s��XżRċ���9ȉ�U�ۗ�#)ُ��Źە��v��=3&N;�+��9D�׼.�D,�#��ꗞ�+�u<sYY\��3,!k,�ǝ\��i��ur�Y�7���ƎI�\�P2�ٷ�2Uھ����M�p2�av�YDDÆ}a$>S�n��qx��N^�����^��;6��b��b.�vD��uݵ��|���b���f5�x�W+��᧰���pt
o�^D�����S�*��Q�z�U�Ɖ��1)�B�(�DODǀ�/`����ȯ;�)�e5��䰢/!�|L�e��+�2��[bT�|������#�E��/o��[=��=p�p�q7��t�L���r��XDD�c�rk0���+ξ�{Ka��2��a�$2�e!�,ś����	~�P�삁%�����r�K�1ӵ �"!i�XI5w��u3�-���N(4��ԤѫW��SD��>z[[�ʮ3;y����CH�*!%m��$;�X�ӫ�܌͇� z�B�t?D�g�,b�{�W��C{#������`  �9޹pHsꤛ1��p�-����asp]�}���m���xx��X�༗T��d�|Y|:�;�$�$�����N�#ӋH�@V����}_`)�1 �q��16�06C�H�1O�X�!=(�޶��5B����f>K�g뷤b�S�5+.�!�dh5i(q QQ�0�*��a0� I	�+m�s��i,�Y�U���=m"��0�%S�� �fc�5k0��5��U������hU�(�V����_~��Q�u�o/W-6`u�Y儘#��#G1����8㌷��C(pbb�R7<�Db�&Vr1G7�"��rO�YJz�#;�cdH�*�3�!��E�
i]�����w<��nXQ��f@%짉f�l�dZ��`-3m�5��P�Vi����RZ[���̈Yꁹ�����Om�HńDJf;��GOgfgts�}�,�i��s:��^:+$�vI���7w�\ݍ.vs.<}U��a$H���3a��Q}�VA�Zo�u��ҙ�C���qDw���s�}~��֤r&�3UM�ZK]r�&��m;�Y;�:�����i�F#�w ��6�{{mVѕ�dTaZ���������Y�Y+��QV����&r{�;� �RO���B�4D&I�6�q�&y�ێ/$!�O�N��׵�6�-ؙ_�[|�̈́K&˕P�� |!W�:�y,�AR��P����u�3jC�Z�Wϲ��s�!�b�_�P��(f7%�TGrh�#�n��B!��圑1, [\b*���[n��q�Mb�QNiy�Ht濨�0�l[��oWՅƄYY����yx�R}�Nz�m~����Q4"PĲ��2U0R�Y�u�g)DP�8s}٥�p(v��L$��a�h)�L�h�����OTC!�0��$��Ң/Y�Ĕ�G0
g5�,~��,��̉n�����ڱ��z�#78�,�:��IQ/i�L��Aafh;*p�!�Y2솒$�J9�^r���Δc�JsZ��޺+'h��I%�NT�
�ʨ��g�v��_Cx"<n��X��YFm���g���g9<W	'*��:�4�S�ɸ�%*�K�o-om��wh#l8 ��;۹�E�Ȁ<�F��d�'zǄv����du�Fc���}�e�^0�'Jb��Ʃ9+�ܼ�g�!GU'��2 �"H����I�%������gR��(��2���RE
�.4����-���\�n،Ѣ�U�p�3
�V�c"8yv±p	�7�O؅WC�j�(�6n�Ȫ[HQ�_�0�	�E����f0Y,��)wѪW�D]�dz�j��if�:��߽H͜��^�6����d&�wq��L0��hމP���7i�ۅ��H�4��Z�)�'*E�$DL8g��egX���U1����D@W6ْ�@3]�<��i�O��1���DZ�Si��A N�b����[H:e	�����@o�e�����|�k��a��N���[g��&��.����gT5��{(�������@>����V��?�r�;$���8�bI�V�6IgbäU?��/&��a��w�}�!���9&�֔�/���2<��Jl�ƍ�Q��B����Q#Q^ϼ�y�fJeHji]Z�7�J��w����/��u�Ѕ}X:!\��n��{�gV�ө9]ސ<ûs�
��wֺ�"%S�o�Z�s�x%;ԇ��	��H�;��b�;T���M�a��y<u���6@%�	s�E���m��<�Y��{���)`�=���k�+���*��aI��Y�H��1��ۼ^�0�.�����T�V�e��|D#4{}�
>�mSf6[Q��f�u��4[���c�T�ܯπ�}��xC���=�º���y��+����MO������36%I�	!�ۖ�m@�M饹����k/�B'�M��-,�^Z��LΣ�W��L`7tK��\ӳT�K;
�W���:�3)�a�o#[A~7ץ�Y�������QE* �%��m��m��(��(�1D#pH�e��&�MEm�
(��R9QEq���$qSb)E��!$�!H�!p���n4�%��Q�wffh�If}�I$�݀�ə�� (.���c�%ܟ�x�������ޒI {�{�W�ӯ��*�8�A�UvzH �H =U�x��|׌�����9�\�2`���d��dL���3r��]W�ڈ���v���Z�\���7i�S��d��aĕ���B��w$ૂn�K����,g�s"|�E]�»V]7�;�)Z����Ą��K��Zt��s�cט:VX��;14�%E�q(��EQ%E��i�#-���B�6LIF�,����L���M��n��$�@ƣ򐘈b��ڄ#,��P��J�ME�e�FD�B4䑟)17lH���!e�ˋ��K@��\iRE��m�ؑ�"2�A��a�-�ӈ�"16�D���K��<�r0�,@�-����2�QHbp��J)�(������w&Z�����-��k���nkBe�����C=�����7m��:]��w��9ҫ�B*5E�F����v5�ի:��P�fW:�	n�]�@�P�5"1>���'y\�ř5�g�-1��qs���5r����wBX�:-@�ga|,�]�2X��˧A���fZ��\�Yr��;�6S]��B�U]ULpG+n�t��K7�����~�&�W����&�Un�Z�I���Be����(��خl�hX(�k�s E�&,gU�u�e�O���o�� ���iƠ �V(�^u�7^��n���K3A:F�����:N![�U�zTkP`ݫ�b��OB�A3bA�l"H�wn�wϽ#=��YNF�����G"bEҺ��:����T�� 1>�T*�=��Dx{�i�F�cO���| ��/TVI�3�;�!�Pd����nn���5� � �{���]L���M�T2�1=�����&+B�p2�LH��	�BX�t�o V�g���G�=J
�ܻ��a�4<[�9��]j�S�:���*0�����3��׻ȑF���Υ�3�N^�%M�!����D�d��H��-���~�T���/D!f���^+.��D�/���{z9���hK�x�L����>�98¡v��?_/_-�"slߝh��g�3@Y�x0�M�I�'7��YI��N�fqg��n@)9{�gVR�F���n�P�3o4��Hm��^z쪩n�!Κ�jJ�I�%����Pr�����\�[�M�"�F2���7�0��x
����*/�BT�C�*��K�C��S6dp�s[1'pH]\Ͳ�a0ٸ.�MK1�΋�uHw�t��y6�8z��jԘG�K5f��Zl�&��G{x��Zū�a��7D�(Q�����z9n�遗B��@�&�h(h�B�]^f�~�sԽ��J���3��O��%&�JH�!�#�"I��Sd.�ى'�����s1�o�e��]ݘ�=YB�X�p� ��1'�HH�&��b1��i&�1�m!1+�s2���+;[��tW]n���/�{�� ���>>r3�#�mvm�g�f�?$��c4k̋��B"f�>0�;�aǘ2���Tl�,�,b����p��4�2�-��d���ˀK�=z�Z�)�����=��-k�)���i"5Y�^�Ω���PWIERX[�u��L<I��ZR�p���v�)N�FfH�����	��qQ�����'��Q �C�L�$��YP	�肅�F��y��o^�W%1��gVR�F�^�[-�)�0$w�����N�:y�*����4jq ��Tj�sQ���H��lh]�ʷ�h`�5[�m�{��q�P���&"����w_{����뀑�1���B!�������k.O�H�`G��D����b�JS��I Fm勽>�x��$Ɓ-�5�v��]��V��!ׇ�W3�r��;�q]��B���Њ�^!�����D%�����M�=��R�w���w&-<G
�(���\#�W�%k7\�q$���	��=���b������
����&��Sy�j�l<�.�܇,4�H�����~�����;qϬ�<�)D#sϤF*<�]_ot�"�N�F�����$Y��a��H{�z��w<5��l#K���\c
!�0̸$��������fzSa�ņ��zd�p�;��=ǆ�9V[�t�	<�
5������CY�W~��Q�$�H�q����(�8��cJ�a�ވ����?��Wb��͡vQ���=�*�Q,������lc\	һ� ��B�Ƞ��mN)4kv(͔��D$I�����{��@��h��;�2�{�u�>Ow��x��:���d��4`�����z�ꬪ���2]��v�2���+*�3����%���+5!N�4�̵���GĂO�xy�Ii���A v��7��W��JRJ���Hw�d��W}oB=0Oq��t�����i���-¨��nt��b�sM�K�C�ԃ5��!nv�D�%���h�n.��ʶb���ꗞF��������^2{F�4V�,�Z-��ܻ�a&��kL�9���nQ��A�2v��9b�%(�nzqo�K�Q\����?7[�+��p���*;�~!�Uu�ő7���
)J\=���VƋ�L���yr	�	x/���ZÇ�N�O�Uq2�C�6�,��#M�-��6���U9���y
9��Ď���c��j��p���l������π�^ڍ�{p�ʯ
���_	s��'�����õ%f-b9t��'��K'{��kDu�1�f��ۇ2���I^ �̨�:�%��A��v� �U�e��ȋhJ�ʆ�Gl9;l/i��5�S���~���Yl�p$jr�Ű��s�kui���"7L��R " �4v��*�8�b��7H���!�(L�����I+s��`�9��k���+Z�E�xJ�ئ��x�D�|NtVŐ��F�p�3)7�X_r_���y��Q���b-�on2���ь��c�_�Nf����]R��ѹ�Q�RauT�i�~��o�ɧ�V7�nՂLe!�$0W6��ԃ*i֫BR�	[dc�w��qB��8��V��=�Ig�C�0��4�2��X�`vLA��v�b�Ey?c~�> ���s��7y�3��j��߉�����HQL! ����N㳪Y�~�]8�ϙ�ffkt���K��T����T��&3$H���4�ED�f!�EG�e�h"(��!�hc�����J�Qnv��b�����q��D���M����وI;-��ۯ��şo϶�"�p�Ӓ��Z�bAm#�@��S�Mfd҆@�	�����Bo=&J�����Cs�zE�;���g^������v�i:SA�R�3����#K�<fѮ��[C�sT��^�+$�v,�I0��VT�}�,��X9C�� 	��3,S�R�xDG59���r�	���.���@�rqo�����y�H;�2SP�j���lh\�*贎�D����8=[�l����*�nK����,�$q��Y�U?���][�{F23U�5����BU��6���dΝ�p��3�hW�ey�(^�zN���iRsr�����˥�Ϯ����C�����͘��u�Z���F-y� ��n9+�b�����H$A��w:ͪ�sR����\�:��Io62�ˮW]UPT�D�j$�P�0�A��j�	"��r��X�j�^�ң2�,��G�h��$���h�pі�h�if��&�OAܪv-P�LY�z$0yBR�k<�e������T`�V��F��&�#HDK�)Ο�s{��xH�Lvc8�&�Z�K�pz{K��%��aW��g �Ң/Y�Ă�HA�C��F>_j"�x��5�؆����I�ԣ7�����y��N��ĆG���%��㉅�S�o��ܨ���+'h�y�0�YY����<00�nΉ�1od"��M1ns��N_�(�')Q�M��6T����Ό�x��A��"�(�"��cJ�J!%���J�	�
;��̔�4ڢ(Vq�8m��<!��BԻ5��\G˂j��ר�E!�@�>>��� ��#�`�k]>���񧛫�N�6^W�����ʏ>������K˒9����W^�/y��{]oxq@���̍DM��������x�w�K�bB�� �1���\����W��$�M�V5Z�����6��7v`ƫ</%�!�
����Z�(B;i�F��Fۋ6֝�,�Z-��xV}�e|��v�-���E^	P���V/����X.�~����%Ө��;�ycHdU]@�1$o�Lyw�GRN�D0@���s�f�غ�RS�
۩fK
#,eC܃;�&�9W<�nu3$�]�&�1k!a���[%�$<ci/�i~�Y��89�$���={�a�N���8{�&?{��p.�9@��F���XۜaP�ɓ5��}�ߟ�֛(p��uD��<}��g��+���`/�W���>Ex�����)܅�b�{���RC���:��m>+���	�o1o%L�����֜ݨ�������]N�޲O03Q�������YLQ^��K}�{�P�Q1�|��W�4wY���t�ѬW��Sĩ�w���D�S�U�Y�IkF�����޼�eU�-���ˠirޓtj�ԃ�6�C�����3:;�æq�)>#[#����i�m��L[1��p�)��7m�vb6���:��P��ld�b#%��gE亥��[��K�ǫ�d�ty���o�i��ٸ���Ç�����K��>�(H`�J�ݍX�b���wٽ��}eSl���IPS�;W��B�^~��H������J�iQ
K�����>��v�0�\��Y(p�ٞ�����R�t�Fe����<�ލ/��z�����0m^�>+�}w�g��_wB�cDE%$� R0H1ƊF9/l[c�~����	$��%��_^V����v���P����@Ph2�-@�n5$~m��M�؂4�b'(�ac�����J�񚂋�2�6k�� ��p��g�4��u�k;�|4�4k�/�7&�$�T7�G;Pv|��w��|+[SM����K�l�HL�o�_�����Tlټ͈�}H� I~^�p�D�,���Q��;;P "
�]�H=�ʧ�q�E�e*iq�Th��u��ԙ�C�޷{�Q���Y;ʹ���4R�ˆ�]�m�f��I	�Z:,VE'oIjA���!WL���ˬ��J/�m�Í>��!T�}��V�k��{ު���m���N9K�9��!�Z���j�eQ����i��7�F]��hQӹ���,��ֿ{�R�u$1E�[I������;T^�y�Q�T��g�/�*��k�nN>���.f��Ô��ICul=��&�N+�RnU�cb6F�N�V��V�D� �>���#2��'�_^�ûzi�=b]�a[[�����Ŕ���놾�XԽǏ�.���D{
��$
m��Fk�o �|^33 �{����A�Pj���S��%*l7y;�a��!�{�<��ǰn���S������e�l�"�_P*���)o㳕�b7�x_� }݀+̒s��˚K*l�2���!X����-BrO'�_'�q܇pyy�ܞOR!�99 |�{Ýh��Mx1@Fs�����t4�x�� Y��c�/�����Mg���#�[�4�.�&����'��$-��b�U���d'Gy�MnZb�)�`�z�P/����,�oO®"7fcp���h��]V,�Ȗ�?V����8�G�Y}L�M�@����xޣ���:�a��!V}V���hdO"�o�>�����<݃Nʛm�Y#�sCYx�&�#�x�=I��a~������Y��%n/fN�^�-�1�y�vR�c��H�Wڗ5�-��?l��)9Q`b32I���&D��A$I$M�.Dr�h��Q�l�m��E�w�����۽$�6낇N�����	&� 32G�$���.�����ɷwv�'���݉wwa���32@������� 32G>����>�N 2���o��y�y}��L��QŃi��vR��m]&K����z�+aV�S�y�@�2v�1���h{y�N��0n`f��.b�i,�_�ݞ,�w\��٫����o��}�t�Zwxe�PSB2�[)�ˍJDUNں8;=�C��q'�9�k��i<R�,��Vnv.���)b�g]�\ޘ�8V�|�܁�	a��(��p��r[$(���Q�I0�1"�m�d��H�
���sɐ\)nB`D��e�j˒'"�-0�M��.&cA�#M��7<c�E��$�Bɂ,�XjH�
Q�I�q���U-5��b��,|�cD�y-�����N�qrᴣ�D�� ��M�ٷ�����ՙݯ�-m4TK��fA�
;u�43%vj�R�pe��kV�e��j��Q������Wa����m�PT)�J<��˲����.X�dʆ�$��]����+�w[�C��u��)��_䗙PA8��:�T��1��8��d]��z���$�g�T^kR`�},Y�u�Ң_}�&$5x�m+}H�7�Ǵ�9�C���a��*Nw�&�#���S�6ũ�t�>�8j8�ץ�I���f�R��ߏ��J2���nD2�T����L��*M>��;/���UC��M(���q4��\���\��-����=~�P��^�b9|6ܺ�{��:���.=r�г��#����5D�R�2�� �u�K��~ �f�2���ʸIRp����3+H�	[��t���n��dx��jFg�o�b��v6�NE�JA�N�+��\�}���{��X�
�[�ZcCO�<���UU��Ƒ2�D�	#e7iI��ؼ�}ה�m��e��1TN�{�a`��}R�(�X,�J��m%�^t�9�\�8�FV:I��i��2�%?�����:0$���-�T0��Pd�k��i=;v nq�$<.�^!�se!u��z_�/ ���'DAyw
-��)���b��K���v]����"8���J��7����i�$�=���jc�r.m��A�c���ŭ�Z�ʎ�u��!A�g�Fi�x�0 �"i�cJ��Ln�:�!2l&E�t��#9�%M��RD;�c�p�UB�ˍ#�~���,U�2q=B��Rd��-�=Sh�*¢[�1��thk]\��ź����29R�\]�b*��Os���i�B�@}A�$Q^���ƛX;��mSWX����gk���$�eܤ�aǹ7��^��|���\B�;�w�� bD�N�:�+�b�TӰ ���A!-����uW��؍庤�
�ܭQ����]�1չ�Y�l�)R��vJ�BL-B�D8�����66����mV����+6�L�T#��k���H��5�jR|�cQ(�r![f��c�3����E`ʇ�W�B�YU�D<�(w�q��(�$>fw<��W�]Q�!�(��Bdn���[�露�2
�MC M;݂��v��31!�*�oIr5��/9=okk�Q��Q�&j�ь�we.��$�Z�+)�x	���u8��cq��ű�Z�Sj��_3hs+�DD�2�*C�D�m�9�X����6�zQܹ0�R|u1����͕]�o���M��Ov��J�>�ӛ�и6�.[&�z��=�q�#���{/�e�w����<�9��Z���d��L��i g7ջ���
2w�el��UB��dtޓtꗻ��	����ǲ����HU�o<�T䷉�yv±Ph>3�n�^S;��a%0��1�T�Ѯ[�~^n2D�T((�@��E�����!�����p������
��ӊ���"h@���ZOv��)�	0|��f�`�J��X�U�6�*�K[#6˼̜�h
�r�p�� �h-������X�2�ЅMՍ���Tt��t��N�s,	�2�Ӳ��DC�-��J�8{ޭ���ۃ�dJ[�!F��C�q~��+�w@���-�-��)�q!���oIu���a0��up`i���v2]��#H�p@>7_����[ �IƊ0��� M���>�l���I�	7n�1�(�d9�_e6���W,lƉQ�Ӊ�\`��6��R��*32�"#'�,X��9�9��Al��9!<��/Ge�H�0��^�T՗��4v�b*�w�˒'�al���澓`'}����iL�N���g��܀$-l��j�Th�,�;-�e��5(�*��5�l�]��"�BgXҭB�BK5���*���
��Z����2~���;�^����ۜ���1|�Н�D<�d��b4�M�=�5�2��U{. <K�؊�a5^�q�i�Tۻ"�8zo��h�ty��9�F\�;��7�K��o�$�f7���ƈA���Z�w���zN�9zPu*{QŶ^nH�mqL�<�w��]�w`�LX"��3�WJ��q!V-���s�C��=�@���T��'��.���w���V��>2��҄�%�����ܙ����ԚS
}]�ˢ�gK���ė�W(��W�@L%H��p�"2H�l1$2�By��HQ).��oe����PH�5�ۮ�����*5F��&�u�2k��-(,]VXGȬY���n��$EH�P�RC�6�Q���}�z�&ȪTk
� ��2��A�Sea�xT�w#gC)S2ޒ��N��aA�&k|=M���Uxi�.�k�����
��7F����y������[2���5kr#4�D(��H�!�*ë�+�r4�г���B$���"�U�߼���r�(Vq��l��hh^bҜ�-�z�|l���i �X��w<��p��@J�]s�,���bZ'�w��VB������%ƝW����w��3��5\��1�i
"
��{ÄE[��s��%-%���ԭ��Q�[���aM�|�>`x�G�e�9�=ï7��뮅hJ����JUn%���14�?=5��k�S��c�N�K#F�)����P}�\�f�y�a�u�˾c�u^T��œ�B�/�KR��õl=�䦤X0]�j�+����&��F�"�d��dݯ���W� �j��b*�\������y$�V�j��֨
�2�kI��gU����mh֡64
���9
"�,z��e��U�<ç�=h��\���mt��< ׌���=�i�W�yNڸ)�����+�O�V�~��0����c��!�NEm㿿~�46c)Q�v�5�]}��h�ͯUi�b�z�șg�
�eN�X��6�v5��xz\�V��f�d�m�9J�b�~�31.`"$�9j�p�{|[g���u
1,U(d�C>3,k�:���/#f���&��/IjNv��B�*t�^��K�<I>>>�8��i7�p��$tW]�{��!���<�/���� ��5�W��n�i4�Xl��c�hV�=��+em���2w��JwV'W����Y�{���@����0|�G��TM'��d
��J�[ȱI�^���)��`0���͆G��ў����ʶb-��eHQQ{[�+��2{������`�*T'6��\��e�����33_�{���D�~Uώ�Bj�5����4�J�2Cl� _��C9ݑ	�o=H2f�	�L��֤��3����-����b��w�E-g�k�(�-c�`�&�ϝ�!����~��^��D(����D4�`��'���|��x:0L��`��G)M�1j�XG �W���9��ee�0�PD̵V2*^�3'q$��T��v�W���� ��#`	�[%j�UO��}9��v����"i��i��z�/�5|~���*��CX�rF�.D�)�qE���U��<�Y6�m��$�V����m��!7W��ɴ��*3�5 �!	Bd���bs��[�@�-��B6�����ٛ��\�brB�}�؇O��P�2
�'y���Eo*�eABv	jnA�)�y�e�G� �le�>T��;j���2�$C�4�ΣJ���c
�P��@�Le:I��߳7��*�4�!�ms�o�d�|�}����`#R@�h$�D�Χ^���?S`"��Q�Q�{���7�dQZz*��js%Ɂ,.]�24nP�'v$���/WkL�Rʐ� ��<��0����~G��2����ah�͛(m-�UR�(�v=?QC��g�������U���$��,��s7	�A�8Cs�b��C[i�JgU��"Z�m��2ηY�ˌv:}eA����3c��3R4e���2nހ�S4S*�%@��	�����I�IB�l+
� ������<0�h>��%R�s'���p�~����x�i$��D�3>ϕyE2�tw�����>�6�}y]�6�eݔ�`D"-DZ�b��Rb��A]��Ք����٭gWV=E �h�{�����2�nu�퓸2k!����ܼ"�^��[���z����,]�1Rr�!�Ps�ZDĆZ��$9�A߽ٶg�s��D�6fUV�*�h�oa$�����v�GhOxՀC��3%��S+d�G,5K����Z\�Z���<e�CD�$��a8�*��ڷ��[�7�GH5k2��mDP�2�u���x�<���'���9y�Em� %��%�Oz�p�X���7SV!��&I`�J����ѳ&F5��Y��J���x���G��l�?�Z}Kr�����2���kx3T��>2�d�\f�E���]e����ϖ���W-��H��.�<�R��Z�Im�u3n���b��;f�Û��X
4}�P�h]�Omi�(�#Ӫ�t#��e��Q]US�SQX��S��ӳ]�r�R�{�W�;�፬�dF��r	FET��ed�!�V��
7�j�*���=�"b�5����4}?5���:B$)�!,�׃��z�L^w%�h*{��bZY���Z
�+%7(w�z���DgM�j�lQ�>�7?�{�h�ȇ�燮��7��N��%��RD�>[�1t��]��6w�!f�W����rBAy$�CeKaX���c(��&��F��(�n}�ᐘ��0,�޴�W��bÇ�N�Q��U�t�Y4#���DY�M�4�kPj�B5p��w.�y�����j"�j���A�a��Z��׸wo��gm
j"W�0��X�T���<6.�bl" �S��M�LY[%�hѣ��R�3��1^�ѵ��#_��p����A�(h;�#�7ňG��p:Ӵȅ�xt�~�b���[Q�ٱ��U��S<K~^�zҙ6Ц���(-�	�E���8��Y��۩�]e�U�ǧ�~ꓧ�u`;3��ű�S�ddza����ֶudԍ^�ǡw��"��y?�`i���8�_w���%z��]�1r<$��s��5$�p<>�ʻp��a�1�O��O�$��>G�e�SN���>S6in׽�W[` σ��o�h7�m?�5>�X><3}�/q^�C�6A=�����7���>�M r����>�g��f���s[c�ùd�ҕe�u��{�Ϫk�P��O8ښke��Ę�&�{ƣ�,ְ�� 'g`�8̧�2m���*��&9��u���>�(�M�Յһ��=yY��xn1"��6K�T�ξ.���Xu�)�9�ݢ��A����4r��9l������ւ��9r÷I^�u�e�uY9�~�C8��H&َG�"�lq$�Q�.EQE���Q6�QB�j(�2EH%QE��QQēI8Ԍ�.'���̒9j��H�p�aH
'�9��Dq�s���� �2@I�����q�
�R�v �&fL�ǽ������3$I =���{��|��U`9�I6���{�@7w` ��T�n�=�'N���g5;�쬻}7�ܗ���On:�H��o�鮮�R��ëM��J��ݡ�i)����);�(gh��rgF̪�5��"�Z��y~y�����p��O8I����w��wD�|1�����*M�׆�>�Rt������un9�WG�k��$��|JMER�5FKbY�2Q)��(��0����f$�h��ϣJ6�)؂1�"�2GG�4�d��m�B���M�ȁ3!���l����P�D�^�#!&FT��Ci2Ĉ��>��P�-"p�˒���XN(�D\-�r4
AqB�A�၂�P��-7H(K�D�$,���P8�r R$�QE+rس{jzƽBd�S�s�����v��ɜn�;��ՓR��}؇v���Z2�y��\xn!�Y�Bro1������)��h�۫�	T�>)e9vk��RJ#jBZ\��o���#X�m���ᨓ]Ӓ��9-�6���)�#�Y�; �q�^R+42�����4,f��0���W6oaM���j�g>��nc3p�]kݢ�/�J�:���o�o	/h�Ev�+%�������N��ޕ�nR^~��x �� 9�-ŋԳ7hOx4z��ـd��A��Έ*�CW��D ���/���ց!s�����ܳ��JE ��t(�
��%&X�P=��0E���]ݷ��8m���F(�J�Y��Hh \��?z��VʳJ�)�P m�̸�RL��qʡf�/��E� �ս�T��DT��TV�6�+	��u̴f^�����34)f�.å�����^_9@��3|</ ��O6|-�P�{�1�h�̴g*�a�m+�tt5�r@�*!�5�*z��b��Kܼ�#1��Z���z���tK��JH�;0����j�.xY�N������[�gU��
_j �A��A�����w������Kʼ�1�]�c�Xz^t�Lu (|>>22;�"'Y�G#\̐�������Mn�� ��N�si�F�9J֝j��Y��V��|f��g,��<< �%}*���ڷ�T2�U���׬�k��������{���EfFHl�30r�] 2�T��}�W����Z.C���QINǇ�=���v�!Io����v�sl
[�E�~@�i)�g�������I/ ��#R�k���v��y��(UaoN�tf!�Cj�t�y ��/��]�r��}K�,�~�|�B�&e��}�&�X'z����L\��S���U��a��dD��\լ�(�6��Q���n��%ᘎ[[����a]lMjjm[(l���XZ�&w��S��2
��$f�z�ި�����]G�a�HRa�1��
7cw,zDk2��fdK�H��$�CQGdއEh6T���EnĢjBK
B������ZR�R1�Sm�j�m���19��+x�=]�N�`��e�� K-��C���0��� B�<fO{uc��?3[�2wϝ�5Z�-Q�9�? �o�v��蜰�����,���8�T�^�ܷ�b1*-��H@Z��\��f�t?t8�F�$�r�Y��GLb^0b^��*�Q�,a{ބlf�?/i��R�f�we�vgMh�º%D)=�z�7w_��I�	��3m�� ������{��E�KnR��fS�� �✸mR|��j~��+ܤF`���Є-j�l2h����p&�-�����=�VŢ��҅ Ɉ��I�IB�FV�ŭ��#!خ+�����eϕ�z}����_/ьIe9��A�&,
Kb�]�>|ip�L(2fUU�*�(f]|��> ʍ�B 	 {�z��{Aȏ �=dn뉩{B��L�Z�S�A�9��/��u�*i[��ܳ��M�6��<�7����Y#�*�8�ȁ��A�F�& ���I�l�1ݷݝp�,���i:1�@��	���CVC�����S�0�z�S�H��|vU�\�41�U�rYm-�j'�@J�����9L�N>�l2R������:%��L�$�j��������P�����J�(�Ϭ��N���fl<d�wN9���\��9~��EX�>4c��k��1'u�M� �tTs�"�rd�rҮ*l2=���ͮ�L� �ƬF
B��V8���mU��6�0YR��YK�!��1�\+�TT���C��!���ڝ3x�%I�Ϳ����%�k,�:��)I%��ҏ12o�=����WF=R���@T��|���8��aX������w		3wkA�Dm��Qp�	Ke\!V���+�R	���>�� H�]{���h�3ےI�&,����\� z�����ߟ�].�:]F����F+nit,vX�!wˍ�)}r�sːz��:�`JX�Xcj�#��E!�&OR�P�
�`�N��O���z%"��k(��M�~��kd�Y0FU��+�����cd��sζ	N�"ӛ�7������Ub�;ޞ������s��g.��aA�2�����gs(<I����3����jz���9�f�O���l����z9ߛ.}���*N���'D���p��!�\^�k^���s�%�"쪹�P/U|�X��,k1:�H;U����Eާ��r)m��^y���X�����jr�-`�ШF[�ag]ѡ�c�	�AK0�WHT6�7\�`�M�F(���ku��tzRkm�jYR}
��V���g)p��EWOt��ek��Su���rJ�RD>��d]�ٻwy���ꡎ��L�� ��*��C�PR��������3"AI���6w[��ܨl�ݽ4;��^y�{�K���W�xad�,g�Wrr5�噚�Hky�fZ�F��4��c$@ļ�*hx��>,e���� RxI,�#e��ch|�g7��v0�\5+>s,혝!,B0��h�1ٙ�l�:E8��f	�t�B)/ ��;��m�0%�3���bfb�3Sv���i�ϚT��h��78�_��<�
����$�IѲ59!�Q�Sx�s2j�XD�>�8~;^�����J
�����%@��b���^I��-�L8�݌�e�h�ax��AL�����Tt��vy��)����%����~au�Mbjn[�9�;�Ja�o��)����BwW:J�B��4��fww��2��WLB*��T䷉���/RZ�G�[�z<XЮ����C�CG�<v�lg[I���F�H�Y
B7+�`�!?A�W6��$�+\�ξ����͑N͛� �7i$p8�$�*D!P��HL��b6�J@RM(H�6⌖ʺw��},��fK7q)�8�i�ĢO��D{�=G*Z^�	�X
�S�Y�$��3��Ѡ�3����^S0N�6���öj�������)F6�J!L��]�9�c��K�ΞÅ��k
ӻ�e� �YM�g\�i%l����}�:��0��Q
H��ʷ	�� 0,�Y�帄8�D"��%���d�hzr�pѠ�vߟU��L���Є*n�l2F�Tt��t��#J�50 �ƙ���H�xl��c�����ۄ�2T�J`��aXW���@2şT��lu�B6ߊ"�y��uH~lwX�� m���)��ghɷ��v��by�2}�ȡ����� ���T�2d��`�C�5#>����OS[_�`�1hݩ�g�E�p-�]��yR|�ǌ�A�'Ï�c-3Ek乬�g\j,�\	&�-&��9{��3+6�������\��T�8�s�v�`������b@����Q�$H��d�b�7�s�C��z[F��2�1��uɿ9��Zǳ��I����2g��a���؞�;�l����;���ֱG<�z��1g����ǜ��ogKՙ�C��*܃p҅⟇���wnu��)�pgE � ��ǒu�$�1�ϝSZ�:�n׆q���*W (�׽�)pn�-o�)����|3�Ϛմ�*P^-��]��;�Ǻ|�N5���_a'�s0ձY�zo{�d��<m0
��I�3�$\z;cI�g90Lfs�±�R�J����vJ$H𩲰�%gk0�V�|S�r������q��;�.����Q�*b1�����;}ú:�ڭ�j��p���m��i�@9�6�~�B�y����#�jj�/ۙ"��@���`G7u�Á;���~����T�󝽶���o�J$���.�9f����%�ݾ=*fBNW1K���N*LZ"����
���C3��l֗��d�8r��3<���<���C���\�dL_H��J�]�W1��^�;�����@y���p�Q-6�Oxl^oFom�%E�Y��3OV�'d�y����Y�a��<��յ���*=�-xL�����J�~y�Uk$qvd��,i�f4�NR,	��f,7�t�?�;���P�����%х��?�e=m��_��Z5���Ŵy��_6�΀���G���Ǿ
2�Q�s���fΫ l��Yɇ�5b�KeDA��!������� {q<�:ig3}�$
n�ɚ������* �ȩS��.�Q.鵤��z�i�:L۰��~�y��^@|^/CxQ�5;ۧ�4�e�D��
F�g}�5��6�k36����p��!S���cS3W:��ؑ��y�n�4RH(�� �>dP�j�vPkF��zU.���4���r~���=/�쥏�]|�V�sl
p�3�\.�a�� -�,;ܨ��1��DJh��5�2������]%e.ٸ��W�NZ�uXҬ�~����TV�,��T���,��������;ST(33Wz�%p�g�9٭�l��A)n�U�/b��Νj"��Rd��T�����;�e]o>�4��0��wD�g"Z�[�ٷź;�x�h3��VO�Ǆ͉�y��⹥����M�?)ҠI���;�ƃX(��<#^S[�` u�m�;��Vҥ�n��{w�K��3ۜ����^��"�p-�MDBƽ�p��N*vf� �#���W��6�xQ>ރ�P��{.��JI�=Mk�RY6��������"l@م�#�8�U����~n��Fwco%�5���}����J�|�&2�."���F�H��C
�&�$�̐�-��l���[̾�T���+
�z�XQZD1"D)6A�A�%@���"=d ��b�-P�[��o��,��6����vgMh�WD�D�#;��*��ߢ����L��Z sȓK9�kȬY SD�!,����(T/s,�&Iv�����ރ�Z�]�a���#������2��sԪ4P�ˀZv��v���~�������uO?1g�-�ݷX\>�m���A�p�����7��Ri�x4U�����!]���Ҕ�󦅺>�m8�.����ϨGty���5+�i2M������nkzY`.]�U>�ћS���;m��&��~Y7c�V��B)��=pr�2o;��ә������׼�+6-�e%�a�CT4H{ج�L���BP�c����>�����V����+]��6I�+#�������ٝ���?S��������1"-	ku�؝���Q8����k���ſ�~����6	������wS�����������Oq�꺅�桞���1�� @��	����6�x׉kC��5:ae����׃��^k>r�B��(�:��#�������JtOp�'�O����J��p'r�Hdd���Α����>d�xIO��TK��}�`VƉZ��փw�c^�L�K�x#Z a�I�4}W_5+Z7'�+��a�����O�(x |F	D6���X@i���+���y�����8jOz�ʃ�7'�n�ȬC��X)�5�x���l����f*Е|��S����-p��&��l���.��C�Q���|=�Vٛ�����Y��{��-���K��X>H^p���؁��D���ܜ�ø�Z=������Yg�VA[,b���,��nߙ�׆Ȭ1U�g5>l�DB�K�>t��c����,7��9�% �HK�2	$$Hb ��HL�HӐĜe��d9"D�L����$�؀�����]�n�o��6UU�G�� M�
 fd�̕ �zn���w�.�wrO����=�y�BI��3?>Uo�  L��IY���m�$ʪ�]պ��������i0w���N.����^�Z�n�z`A�Z��\L�pÓ��p�ʉ���3���EKwQ���#����L����o:���R�ɛ��3N�o�f�DDf�C�܊��#	�%�.r�.L`����6��wq6��_v���!�/�F��ޖ�30h�uv$M��Т{��Ԝ�'.[m�
)��19E�	L#!����^�a�rx��%�㈔��I��`���ȨA�H�H�-8Y)�m��D��e��$J7M���C!l�#aN��⪻]�)Δ�+�|�L*/��L^�����J�v�*Ʃ�u6:�q��݉8gc��Y�xA}ݱ�G(X�r��;����xɭ�,^�s9k�f��;������e6�IS����0�(��`�ǻH:������h\�u	����|SWOzb7E�T��|8�.qxWB�G�H��5v/�u����p4�̓Z��;B�Ԋ�f���}%˒�?)�f�O�V�v���i�.�[�s8�b"괩�O2*WEa-�x]�[�"37E9ܪ�Z=U����T���#��ЉI����[��r4v��'���Tv��Z�3f�d��4�6��6�=ǛA��wB�KK�D�v��fi��&j�/�>v�Q�QW*仴Hk�̃�z=�6iBx+j����}���UU?`7n���'�#�����Ne.���خN
��^��%u�薃�k�¤�W6��"ލͺ\�<(O_+WV��aKl!��@ �
�ԝ =G���e���}���iֺ'�|�W�'�
��2)�18��tʉ�Ͱ*̩[v!�1��;�!|��C�\8]�z>P��)��o��rfK�ӭ(�^p�}��s��˦�<�gE����4�P)b#A(a�`eD�O!o�nX���wZZt�A���|R��m2Bm���@	qYI���sZ�Q�0��1��s2+,��#Zs+30�vl�z�- �B'Ă��!�(!j�w��֙	���q��jrO��7<KT�e�859�jm�Kg��P���`�Z�,R�r�zwbI��܅�2*�Q��gXQ�rm��K��z�|��Zp�b7ߔJ�+���n�P}:�!p4��V��i�Y���=Jr$���J���=����]�!��2<%}��,������^w	2l�g�iͶꄝk��&�O��k3��*Hr}�3��X�(a7]&t�C.t?��F~�c���y[��=*�س��)��-R�6��!�߼;6��nw��U�kػM%�����D��&ѭ�Q���Y���+���^*|`}�UJ�֘%�^wZ�	d
Կ�[�}`��/D
�oż�͓8���f�.�4�łgm�{LQ	�Rv�V�S����F�̘�9��PddTE$C
$эKH� @��"Y)�J%��(��`�wA>_�i����4�&��{�l�*��x{�c��W��gG*�2�������k�����v�czw��-{fij���/V�#]K��xc�
�w����['���4T�e��S�Zއ2	;u*�P��ݓ����T��e�J�wrws�ma�K��dk]~���"�d���8�;9w��6ԻԸ�[��m�يD;�z!���ۋ(�j�d[^�&�s<�q��y�<��xM��yZ+��j�7���q\ܦ����0�L����b�{c�:/;��%����>J�e��Y��ʏaS}��|���2K�� >�$���>`��g��	�e:B=�hQ�A����e���U���	�A*�m^-=MEu#�+&i��gI1�:���{g�{�s!���Q�^�k���A�2�!�Jk���Zլ��Ya�E�f,��0��y�Pa�a$VfAExB�>$Ә�w��-c+7S�C�[��d�r�Ꝅ�����9�����/�J�dM�$�}�˯�l�t���Y��C��ǜ8�Dp���	�xȪLJh�&�ٖ������_;�ɜ�d�KtLp��y6^Ad�*$��Y��\��S\��[ w��u1������)����^'�3������O�g83��j�Vl�bZ���\6��bycQfӂe�6M�W��������?޻���a��vӊ4�M�'���%ᬁ6뇫7���߭���lU��M,�a����~�dz#u�SP���!�� |A����|��^5w�5������ЉG$m�\�z'����$ҍ��s*�_+��ĘM�I"��ظM�7(m�)bi� FF�Q)��r ��$眈Yp)A�H$ぃ��^e��S�^op縅2�y�<$�L�@��m�yQ�"9��af�f�E��'�͹a��(;�Th�|њ�1�A��A�	��(�!����q��( �Qb�U����r:�V�%�֟^8��#pG9Y��g�*G"�������9v����s?t�V�K���xS@4
�{����f�ɉ��a�]3D|����}b�;��d����&i�¢��#������7���Zr�;�x�$=qw|T�!Lֿ�SO�};��L�"�=;PƢ %{�=�Ɖ�սȜ�I���U5�mN�Lb?����x��~�Mm5�m}����3g{�7���o�\w@͗J.M',i�&4���1�;�]�s!2l&��g��#�`��k�N:IVcm*�q�җ�]�ݴ���{2}t0�"n�l��܊�*�E����!���;���sR�r�yi�vTa�z���M�MLD�� F���"0bf1i�$ay"�@�#��]�k7�^��C�9UR����q��,l�5��Q�e�f\3Zp�01���3,�̢�Ȭ,����5U�=��1�"�̥�,�h��BJD!i��$ P%%�ط�Ґ�O��]�.\� ���+���Uq�z2�I��{���ku9�i��z����S��M��&'�W���ʺH��yt�Y��m�r�a��{n�7����(䕲ӓ�" '}i0e޶���}��va�*R���u���9�`7l[?\��{��v���fg��R�@S��SĖxZ���볻�Iڠ+,�n��}��6}��e�o{ŉ���P�+zX�`�)651��hV���m�i9���xw?}E��`%K&	$Lgׂ�~���y��j�$��g)���֗Kh�uU5ka�N�y�bv�{�y�D�mt1�vrO�)���>�H�>�\A�OvN3�.%��G�9U��&����nNf*����it�܌rP��Zv��k.�dcdeffcFEY�a����8֓����Q���F�e��"�fQ՛�͇-��
 �0��0˚~$e��I]FH/yoJ�כߔkL��Q�!k�f�q:�����xTCEu/9E�~��,�1�ެk��1'5�Z-#N���[J����&u6%w��{�����ecM`h�-$B�}�a�׍�c>Ȁ�[�;�,�H�%iƕ�xT?��u	����6���&�sp�і�@�xf������F��9$Q6��Mq��./��������z�d�L�Â��X4jLݜ�t�U��L\Υf�Y�;�^�n7s�=�LT�3(�M�Z����~����-�;S��i	�r��Ɩ��׌�C��.��7��Y�����q1��o�z/��7�� O��pf����6�����y���p_<Ѣ�cI��2qx0���=V�UJ���u}9a�@������D @��!F�4ߘ���و�b׉%��>^d��D2��Bo�L��M�)0g�ő���;�~4�-}R�ݚ{o�I�_�}߿=c^�5kg*2M���xfWOC���s���L�D�g"Z�X��M}ؽ��H3;�,�/j�\5=��V�=νV\�������.�u7d;�:|�%\���,u�.4�@4�+vZ3���JسΒ��SJ���%�<��Ob�(���o�[��]�$6�&�!c^N��L���U�׵�Ճ�	����{����*��}t��\�����1��NP�
�9��-�����o{p��	Ƴҳ]�!���"��wZ�'�"8��� < >���p���m�8��'�$6ԅ��~M�AH%	��U]ף#�廦I+#m���wY�/��;r�*�n��LȊ	@\!�zy��a���BƄf6�)��N�r�e�=&LMαiR���n�(�-�gĄ�A$h��$���L4��e@�@�z��T� JD���e�$ ���8d�.6�I6c�TB�������`��ݴ'wҸ��q�%p����[�T�rf
N̙ݕ��x7/��*˪C�_hXZ�pu/�󪈡c�Q�A�۶���������-��H{���v��n��zK:�U5�a\X�e3��Ht�8�\ ���1��+#BSx�d�gI��eU:1�9���9H���,��'���yYMp�{�'7�s�N�9��N���?N�Qq�vb�M&<�V�Ɖ���.&x��-0
͖�D����I%��<�E����.�)�\��1���-N�&"^�J�י���M�B�~�aF�ɷ���֚�Y��qo<ׂ��Q 7� ����A�>���=�(t��6G)18D9*r}�5Uux��Ka������t�Ͼ1������3�uR�F��#R\i�
���p��»v����K�3� �=����'I��&a�$A$-&�-HRs�&�dS>��bvŪd:TLH�&�j�A����T�]i�[*2:�W��ܮ�����U[�:�g�'n�{ͥ�� �sީ�g�U�'ce�őqDL��CF���<4��y�d�L�A��m�M�]U��<;����
gb`��Z��ժh�ϲ�T�z���
]��J�fU:Z!�l�����wg�Y�g�oN^�Wl�b�O����,ύ,�m��Ʃ��x !��[�豭�T<�Q�ٕ�����͹Ϋ{V
gt����{��Zʶ�$�|1�USX��t蘱�]\o6sת5������<E�C���"k�CY�o{�RB28�}U�#y�������i�&lS�!��4~4v!Ѹ�9A$�V�,�dU�uә�b�my��&�Yr���a��7���n����=�^���a��@zQ;(5��4-��TEF]?)�n�����ր�"�1 �1�` �eXA4����SAߣ#��Vf���L�ӘVCd�F�*��Ω����E=37l� �V%�T��i�E�yu�k|�<�����;��ٮ��/L\�]7z�N����˶�.5�]���Ե�����7�VNx
�h�Uٮ�����d]I3�I��K`�fg1�8Y1I�}�Û2��$����y��wB��ݞ��� �-Q|�|=lI?%��+uA͵�6_Y�#�uTb�����
��a���N�!�&٫Sg�&�l��Kt<ʒ,�>���S5���s߇�K�*��ܼ����9��
�uS�j����U]���7td�����͍ ��!�}º��۠cV4-d�qͮ�{Z�T�[��H�y彷}3�y�~;�s7mI�soaޚ�זIV@�Υ���Z��a�ӛ���hI{m׾��Rg�c��gye�lݭѩo:;�Q�=SΧ��9ҎC��|"t����{9��6��vȝ����`>��
e��[����d�g�`[-z��]=��T�0u�_� �{�͏�` )>N���.��8�%�d[k��w�z��o�hy��/�u�����	�������lMU洃ʀ7�u@�r� v��~E����!ܱ���\�NN�\�G������+��^���i��Σ���rJ(.tY�fc��D�J)n���C���B���V'(dtɶ��K ����2�����69qX�ςw�J��G�U�>��|�zkn؞ɷ��/y,��8��Ԣ��zs��+$G������Y0Sٛ�=���F��AY`ث�Q�9r�C��
��9�k������H��ך�EH#LG
EP���.���m�Q@��(�$Ha�G�Y�F�151@��!Q$�-��dȢ�ƒ5)
1��j(�1����f$,��&HJ��w�\u�f��d� |�� I$fL��� ��w۰ �������33�� {�@I$rWٝ�e�2쪰�l'{w`\�N�w` �����ޟH �(1��]^C�Е�wUmCD5mn��Ʊ^b�N�v[sy�����Sg!ֆ=�G-�䆻���n2��ß Nɥ��i�S�k�q��?�ϗ�TY��̒en���>'>�4�pe�f��s[�'�ma�F�ꏌ�-��tim�}e�jӢ�qEQEN@�lB�I5��e�ؐĔ�##�3ID�j8 �@�0$c��P�1��I ��[P2ZRF�$��#!r�Q�D�9$�������!�lH�a�!p"�jB�a��&&��"c)F4R! �"mYm��m�'�F��B�ˊ�9 �L8�(5	i�R��QEH�RIE�a�=�h\�r���\�g*�^,��F����Dv4�]���&�#��4�l��%�JS��s���Wo��(GF�y��+/mC���s���k�D]��ڥJ�����'f��:� ��w#�Ů�c����2�Z3J{d����5��M�<Y����C@{���V�����>��Wr/���;�V����
W30b$�����U:>�gQqn�����j�q���� /D+��A�s=�+��ٙ��E�P�Z��(�#Tx]9��Y  {)4\GNK�+G,�Ӧ�4
�c�C�:��}��f���4- ����x�Bku�6U[@��:[��V�`��zs���vh;�1���DD�R#c�E�����v����+�7HMF�mt���˩B��9$Y���l9wf�^�)HN|�Uu��q�g"6�AØj�ɚ[p�Z�#܃��L*�UQ���]p��Y�Q�V9T:���� x]5�J���-ө�l-ګ�N֜|��}����d8�kr1���f+�W-P��t��Q��{F셴�ntjf�R3*j˖���Ǖf6u����g*�ݷt��μ��7g3e�a"&�����6\RAQFq�(QD�PA��F|��q#;�~����Q����A-�P���3���F�MsW-peF��͝�7힇�cs��J�y���L�h}���|b�/q̠9�Eؗr��3��9��	VK�$F94يuS��u��ʿ"]����I,-�d�x�j��Bɾ�I��V׻�!��*��s��a�93���e�[�/W�٤��������vf�wR�϶�)��F*o��8A(-T��/����������ص�[�k{eNA5�o�L+jˀaK�}x����v��.m��r�����3DRh�&8x=U?�������>G%�@j�~��Pe�hHRRI	#�-��JI/q��ҏ�|۝0�
��.m�ب����)�V�t�/.�ak1� ���mȆ4�"%$ 6�qA!��i�<R(�,�˭�S��s��
�-ݝq��4/2�~���5NSU�\��	V)�h3�{�P���{��=��,5�ZM��<lũ�MR�6�����t5%
�ˢ�����?~P��d��*�w�4-��� �%���.J�b��8E �=�mYz"W��d����y���)���UM������Bg�#a����kf����f���{:�X])��m���g�bX�Y��:b�M&!��.t�M1���[�����=J����}�����ob݆�?z��ns���a�S
�p>�&�![nkU.�]ܞ� lre��ry���-�-E�h�h#83ð\Vfw:��fLW�X�� ��ĝ���ڲ���Y=\�,�tvGk�xu��`Q� x�H�}�c��-9�N��}(� Z�u�����@p���RR0��e^���F�-<�K��S��=���ܥWOV��v��1@�g�i������Q�ׅm�U�����
��|v�h�f������Z��Bb�Q�jIulK�f�
��/��S��(R5{�!o��� ���_��UH׳,i�}��@��4x9s	�p��l�SW���҃D!�m���[/F��ښ�wg�Y�g�Ʃ�-��+���7����{�WE�{&�6���a�BΪW��Ta����Kwh��.�j2J�)���ޖ_����mkF��11,C��oz���:	��uR�]Zl Bb�߿;��cgb�Ju�m_�3�o;4�d�����'I�D��z����~�����w@��l��OO��{��6J��z4&1��&��/*�v��� ��A>@^��6ϳ�^䇆�F%�v,i�iC�:�3ٛ��ՙV5�n���=�K]��N����Ch6#7b��Z��x�F�ITC��(�X����'ȃ�A$��J�NÛ�_�=�����p��-�UR�M�dR�ޫ�{ɣ1=LX�6��z"̷Dw���?��7z`x\��M\�j�Z ��k%t�<��]���V���5��m��E�c2e�7o-k3�w����l*��0trg�p��:�챷�����D˄0�,�^���w��DRh�2�冢s-:�Y�_^���%-���ֽ�7�oST��|�$=�f|n������D+�װ��;.���:ٖ��n}��r�<:sf*2J�)��NUOxtLu����T5�%�&�9��8��K\�֭�ᬎL8��
�
C�}� ��l��1KÎ�l%B;53n��޿������f�8�xb�=�yѥ�#��H����_U�[����U�%��E�BH8�,"��_���\UW�2��gu}��ګn��l)�2?yF�cc���Z3���4� ��h½�ީ�-o �K�e��~欖��k���F4��'c����
���;�C=�{�I���+��UHS�6����:�]��4mCd�d��Y��M�'a�:���3g]��JgS�l�����WU4A*��Kl��K�+�"d;>!ޛȜnS~-Q��̦����4�=�׽��<%'����-a5��qZ8=�ץ�=�Q��u:�;Wݡ�I�ԕ�_]~��9`='Wl��+U�7���EY�0gW�(�}���{����l�F�D K�8�?W�̮p�LI��D�\�� L�m$���WH6Q�&���Y9Q<��z3t�9�9V�
M�jf� F�1j(�"''<g���d�E�[E���v�;�]��P���l�k13�a��g�<<F�/2FmPj��=W}�\����R�[8-�������vq�ExÀC+~ޚ�1`��]S�����$�r��nUT�-;:%��2�d����v�L�Dt4�15����V��:!L�.�yl�uP���R\��*X���"�6�/���Ll��^Cl��pq���ކ7ȩ�W�t��cKw!��(��Չ�i7 &csC�{��']2�HS�6��;8�S��|=�=�{~�m���S�4�6���)�KW>Z����55�p~�J�����ط��V~�ǗB:�.�!�.]�����P�%xML��9<�W�4�ח�k� =��yx@�ZD/?G��lN��+7'k�&��	N���U�׷��Ew����j�����n�t=�26J&Q��	i���d�b>p�P�(��(�B���a�@��D�wk urR��Ƣ��{Ñ��yl��y��Zz�]e���r/��N�D��s	�|���6r��pm앙� �QL��[�ԎZ/��zy��W��=u����.D)����S[����aBy��+��֮l��]���������XѺtLLK�<<�{�X݄F=�u�5����TjN�g��v��4�;l�[ᑬ�3t]AO�S���~��s:w�1�'�t�n� ���`��k���Jˌ}4&-��&8����r)u��^y���`-˂��*"�kFQi�+�n���ni�:�ۓ�݉�j����VJ��̰;�_�Z��N�C����ؐ1l��T�w6�.#"!��r3�j-�d�|zv����T���t�%��]>Ɠ�eƅn7���xy5� G�Vy��Yo;�HfaNV�y+��op��#*��D�8����Y|�<5�7�z��V��N�w��2nXLϭ&�Ũn�9[$ׇ�N6@֮�����e R`�nt͞���c�Cm�é3>�z�R�.r�Ė�C|1��-n�{��!��:K�I@_�s�,���l��K;>��a��Is.�g����a��5�UJ�6hY��T� ��`��E'L�z"Pu�-���H����%�ʧzZ�G�U*�ꢭk�[tKC�r#^�up[������*5�[���2�k�nܫ�g�xy�0�9����h~����L�y[��@c�/B�"�0Gu82��:�G�஥=��c� |4h��^}�wzs�>��}�é��e9|�uzV�L�N.�����)k&�����Z9ǥ���O���26��f��EZ�	�e]B���-6W��U������%�����~�S�v��p��L�����єZa�۪�rz�f���0M<�G=�s0�U�f[�;��W�>R�m��T"-B�r`����F�8���ڳ���N`��n"E�_v���j�Ɂ<=�y+����!;�I�/�j̙n���Z/�ݜ�t�Һ�p^4�9�6j�4Gx}����8�T�OC2���e���c��6N� �6�!�&-��4̱m��]���Ѿ���5Ygynu�n�¸���1v����n�5���'T=ry"�~4d�k��]ft�fmtd�}��,j�d/ "z9����x}G}�0W1X��������1ꪾ� �c+��A2�n�/D\b$���U�v�j/�sz���e����I|�a�H(��y/A$��<D&5�,FdJC
2�~l�e�1��r$�JEU/]��$�	ݕ�n0�����y�(�R�2�;`y��N�L��"I4��uQ_�x��*\�^^��	��(��=�>�s��7f���S&l!1I�)ը�u�Sި���2�h�j�G.��71a��W�B|�O���S��X+=�˞	�h_���z�(ֿg���<b�B:M��.�qtb-w��6�v9w�")�16�&�Ab�֪B�ɷ�"뫯j+=���i��v�y����"Zݜ|wn��S��15�m��U���i@�>�g8�|��= D'�F�{�P�fSDl���s�M�w_"�>�t����˜sV:��Z����<����*����j�����Si3Ė�B�]$�۷���� ������o��0o�`" j�� �����{�X��&�k9�����mPC	E2AWP��"���A\��i������M ���QA2�+J ;�QR��]kDD�G� ��b��Ҫ��"4*��u�a��yu��L���DeT!_ϓ��/�����?�3��������������ϯ�=nO�㑮����?�����tM�.W��������ϟ4g���?�i�g�����N��?���(���������J���B%@ �O��������Y�Z�?���W��~߷��~�����w�T���i�����������u��6�p��&��ӯ�|�W��������_�K�C�'�a��}�s�����'B_�|?=���o����g�����ן�0y�DA��,�BA"��$�@LHP��%!0�BP�!$��	�,��BA	$$�BA	$���$�$�	
@@��,��	�H��(BH���	�@���$!+	@J�$�$�����0BC	2�	$BR�BA	$�	HD$���R,BP�BD�	0�$BL��@BA�2!�BB@A	)! BI!!!$�	�A	$�BK	��	2B@BHK)	#	!	,���$�$�	 @H���HBHHI!$$��H@@�HBJ�JJB�J�B������BB@�J�@���J��$!
HJ2�$�BJ��BJ�!�$��HJ,$�2�H@��0� BH	*2�@B�$�BH��$�$$!*�B��2BI	�HI!$BD�0HD$2(A	2�D$BI)0	$$0�K	$B@BC,�$2H@HI!$�A0�!�HJHH�L��BP�!�J"�$\!)!Z@�(V��J�
B�!��	! ����(I��$������(
Ba(����"X �&����(�"F���"�����*�	�� ��i��V$	�@�F�(����bD&��"&��(h�����$���D������
h
�����)(J

()�(b )	i��"�!�)((����
ZB���hh()*���&�b�bB"$d�H��"�B����������((��" �!�&@(�@�F� �!R!E�%!Eʕ% �"P"@(B�	�(B�`!�aP$U�!�D YQeP�!a	@�� H�!	@��	�%VF aP%@�X�R ��aD�	@�$BF ��BBA!$�`D�P��Q�DaBPd�D� HU BTBAR @`BQ$�$B?� `�! B��@0�*�)
%
1 D!�	CD$�H��$! D�$�I P��!H����+!D!
@����*!,!*,�BH! D���!H(1R( P*@�P�B�*4 R�K@� ��J���dV �@�BBd�!
J�B%BB	@� a BTd	 ��&��(	 �B! �
E�DQ%d B�"�hBa��R�F���$�%� �! 	P!	@��!P�QB�(P(Eb@�
@�
��(B�(��"AJ@��
V�
Ph�
P�
����(H$
��Hd  $HHD`` �XH��HBU��III	$"! ��)!"B��(I�hR��
`H�!Z��JU)T��F�B��f�I$&BHHa $!a HA $T��BDI@$!VBU��a$a!  a a$$$��BHI!$d%������	 "Id!��H��I !�� ��$%! %$!!	R��$%! `$HIIY�� eH�D��!!HRB ��! IHH		HXHI	d!!%��BXIa $$������$!��H! !$!$�IHI	`!!%��FRB��a$Bd!V@e% %XHBP����BRY	����YL�0�K��Ͽ���o���7�������'�����v�W��������:�?���}���]�b~ݟ�����U��z�"  �ϼ�������ø�a����ϱ?����v~,���'��g���q��?��~�����?O������	��?�T}~��W�?y�~��������  ��o��
O���a�����7��G�?�|?߼~�b� ~� ��~���iLه`�g\E@@��v����g����������� tl���3�>ߞ��=�3?��΃�_~�M�����+��A����t������15�'����:;Gi��P@@
-6~���?h��~�~��;?E �g蟵���������@������������?���O�9�������~�����~I��Ϥ��O����^���8�����k���~a������	���ؐ~�����O���O�����E�:>���bI�ž�矷���������>�z$����������|���п���t$OO��`�������|P@@�>�)�A�ϱp_Ow���4g�>��ﾾ�<b���:�����_��0�}{��K�������������L�����3��y�������������7��m���p�����F�_����������G�O���J������}�?�����)��ý|��/�9(�����o����0폀|���؄ن� �� 	 .�@m�f5%U�R6fؐ� "��&�-���   R�6�eYv3�l     � �=e Q� ���5�E
JKZ�JR�HT!R"T�EJ�B�e�"�P�REHP�"U'�jRKZ(��	)T*�*m���R�Q��)m�mcY%Rm��j��T�ϔE�@��Ѧ��E�t7+j���H}�=e'��ك�u���Uwu���;CgnP����wSn��Ɉ�I�� uQA*�K��p P ޸8   h��p  4�� ��L�۝��'ep.�V��ہ�*���ԩJwKr������Ԋ
�;�>�%H�UAGx�nw���:T��P${l��iW��V�=;קJ�v���u�.�iZ뇻ޏl)���4+mq�ҭi�:��I��3�@�P{of
�*��`]��u���1ٹ�X�:�v�û��:t�2�]��@ژ ��۝ٻ3u��T������@�T�){xlws�+�L �A!��
Z��7u��S��t5��w �5L[����QP/���Y� ��7z���7�����ҳ-lm���@��Q�Zΰ��D��1G!��wt��V6Ν�_ t�@UP x�q`�6���wn� ���������@�\�@t3sp+���(Օ�sS�sx:J���4Y惣��t�˷uFA�����m�3Q��kY`w_pi��4 .팲I"> eID (U/��@�H[�NV tj�� �{���Ys8n7F��� ���rC�.n9�A�8��r����Q>�T� ��{k���AӀ��t� �`��$��5� 4�ӹ�N�]ոh���h                 S�J�        ��1�Q        �M���UR�  &&	��d�LO��h�4h!�������?�%U        	5	R�h�� D��d�Q��F�z'�?�������v��G��s�dL�����E�Ww�j�L�@ ]�����?���@�䒈��HH� ����?���@ �d���������/���,��9������������O�Q��y�&?f:��~�� � ��1X��W?g��� ����*���P~V~8��#���X� 0������]]~��'���~�� @ ����҅��Շ���~��Z��ۻ��K���]|��4���}��ۮ[gk+����O���z�-��s��� R:ӷ���EO\O�٢�)YN��2����5s�g �i3���d��9S�:�h�c�2x��N�$l#��[zK�ߛ���elۣ���o	��QAN�gQ���CV�ljtK;% 	�;.��Ǘ+}�')�y�k��i�_+e�2]��XPU�"x����r3���.�b�U���E����9	E"q*�	1���Ըͩʬ��'��yis�μ��ɺcU���]ǳ$|�@������1K��FC��D�+��"-Sg/M��墖,��.
h��ͶI���B+Z�E�7re_Ğ�zp���Mn�ʴ}K�&�e��fj8�F��Z���E-t�%QL]j����:�q�e�R�R�9SQ{V���-��'n=�׌)iY,P����'��="64��F����OH��2�QzN�}�cX��i4t�n�K3(�u��Ḁ�-�rw�c�����y�-I��_<�))jѾ�K�u�yI�k�<�tyۯ��^c�d�M��"��f�~��/1�w|�ȩթ�Qֵ�{�Z��8I�9�����(��5���G���E�X�̬=1�TaW�:�M��7���P�L����V��Ȏc&:��Q�s�=y^6I��v�$jԶ�J��Z��L-x�����kGw��)�����.V�&~H������c�w��UST�{��1UuH�ynϩݫs_X_6*�*g�ȡ��Z��G�Z�N<:딗��9��'�[���^�+��'�c]h�xn�E�K�V�J����0c�:zr�1�vbe�-��ձ��M�0�e0蕢͍6P^��T���}�b9��Dw�<�� �j��H���iH$��Iu/8����R�ZƢ:�R�1N쫵\�9/9�����H������ڜ:�1�X�J�o�����ϒG3�Hࣅ�{&ѩBA5�tZ+%]i̍�GTv�(�Q���1i�����D{&5� �˽��)�%�c�V��Z1�RK�1NX����-=|�Ϙ��ɉ[]K���R��Z�>=Uj�D���ۗ\��5O�u�Vof<����]m�j�g�umK\;ݮyIպ�ɤ��))��.�	Gy�}ߪ�����]G����,T[�ʱ#�K��ڏ�SXĥ��
[έޥ���%��]m�TL�,R��%�u�Z�����v�.O5�����-�VLE(|%��=G:��T����:�lc�w}\��պ��EDj]J��s�-)G]�JX��+�ok��ǅ��Oз���L%T�}�z"�6aⅯY�%݋:m�0��
�:�D�P���k�8��ڴ�ݑ��-��<����Dݺ5I�מ�S���/��y���m�j\���Q{���ξ�W�.�"�Ҙ�{GR��twu�Sd��ļ�5�[o�i['Y�����D�)v{^c��̭,mW�x�^y/��5[ y�wj�n�κ0��SUz����xy�RD\d�i-c����<)�\���[��V�bj"��D��p�e:��C��</(!�:��j��w��A�Ẽ</v��\x��.ㄟY&�V�N�Z��&u/\d5+sͮԭry�=�v��O��Ssc��y�C�Ze/v��S�Gw��js�<�W���{ʣ�m�RRJ�_V�)��y�9�Ȧ猪���[V�ך�ߏ7}R�X�]W^�%�Q���v|����D��hյ����-֭Z�+�k:_������t�܏5ȵ��Uu)x�4���۲��
b�-�Zx���>N �%)�8JR$� �Hp�"R	r@ �)��	 %�ĩ"D�J@HD��"@�*HG	 �9* J\A��|�O'���zv::�c�����+�ɢ�>�b�#5E�$���) ��b�ǎ�l�U^v�}��9���r���1��|���q=����a.�d���g�a8IcMЕiER�ώ��BNQ"a� �:h���QӐT6`t�>	u1��П��X�F��>j;|�r��-�z��K7w;|pf�3�>Ӈ8aӺp�ȅ�x{ۜ��WM!�4K]��R���)ot����C�_����u���ZT�k@uo
��T�Vm���n䏊��a��:{Yj��t��
�NF4�[�{e��E2"����eA��>ס�mŚ�C�Vu߱-��-qmֵ��-� ɬd�J��--�/%jַ6cҞek��5�5"W��E#�1�;[D�v�e�.��sh(�-oF��"�v��YY�keFՇ\B9,֠�;�S�܆���m�I_R�Տ#��k��y�-ћik;X��	=fJ��ok5&���Uz�Q���9P�3THg��h!�^h!���b��;!�:���B$#7h�l2�ܷ��"�� ���{R��um�BΠ�v՚ܘ�jf���d�/5��0�z�c<�ٲۂ���䄪ܻGmV��f���&�o�LD�-�P�B9l�H=OV̅˳aY�47��dOU��%o*�2��6����7���
��zB��ֻt�fH��LC��K����D��k�A��Q�;�+Y���+M�ڋ�J��:J�tւnfbn�5^
�ө�8%=�֖�nkԶc%1{2Y;f��c=����o�i&X��,����w�s��}�wC����h�tC���I8���4�n���x'5�כs3"4:i�������")	e[����Yӯt'R��;,d�0K�R.���Z��ż�jES� �\��ԋ/]������kiX�E�&��5R�wq��RKr��*��Zw��TF^̍����A�#�1i��S/�Ɏ�\B�����U/��� � 5W��ۛ�Z÷[@�D�:�i���^�����=h��]��\珇'&��#w�����56����ɴ�K�W�W�e�]@��I|��xT��]���e]��hުAėM���o^���۸ lܔF!q��r�\��ڽ����BƮv�;WSo�cg98*�mJg���c����L`r������K�Hk�^qa�N1j�t_3����e�.��~�&m_'��]�������<M���������AD﹋Է���5� ��:��i���u�Q�N�1�����O;M�c(�:��9b�9 W�o����=��(�1[�R�S�ɷ�
��o�� ��n�9A��ۢ2��Э��1��r��{,@������6�]udbƴm���� q�Wy�19��(�V�l��z��B�q�������#���[N�^��Z�:h̎���O.I��&'�r�0e����tMfT��1��BKE��L貀{����$ĺ`p%zn�+U��;xuf�"黗����CX�T�tha�;�K`X�T��7�LH�nT�68o��n�fh��F!B���2����;��٭��\��oy>��'Tד]*�����]�lF��$�:��y�*�v�X=�xG�UL�����n�XW�{,c�jPiF�
B�����z��!P�b��	bn�N	��ˠ��~�*�l>jؼ�/�Z��)*��6-�ع�(�4���k��Û�S.�^��͙7-j{P68sr��ñ�LW�X���e�ъk�*R���t��ioj��wE�N�&&���\�!��xfMYgPö�p���U��1MLɋ3��@/Bk6�l3]b�ܨ��m�6���X���){����םX�L�n��G:K�L��� *�b}�:�/8<�]��2�ʕz��ڻs�2q�ؑWk<`�;��%]��1ctlXaM*�
�9�_`�a3��m�X��<aPټ�[V6v^���ڀ�4<*!�V���< V��/J˖�Cʪ��)5w��c�g��l�HJY{|��u�ګ��먵"Ɔ4�ۚƗ"���`L�+���S�I����l�A��n�����wyL�e�p������8$d�7��I�<h���ńb�e�S����Uvl�T<.P�@�sW.ݝ����ue+ߪh["UB�b��M��}�v膻D1� �V��P��`����vi��+D9�Ƶv��,���S���,����TC٥��r��u�0)Y��%ܣp�I��IR��e�Qk)evǣDD�勻��Z�[!�6��H�2�"S�깛)�7A��[\$���EY3��M\���R�d\�K��L���d;�"�Q,5�Gv5�T0*�ݴ���7C��D3�!�����+�yӼ{�^2����T�.u��tf��
\13����e1T�����oiBY��6��M���$:$5�!�	����(�n�lHo4B�D0$9�	�T��D+TCbB�D+4B�D*�j�7A1�!���C���]��Tu��{�m�=˔����8O�<j�����z%��uZ��
S3'Fa2�,�GK:�񫔼Ǯ�_�ܵ�˽c�J���n�*u���EGS�S�
�k��1�sWӵ��T�1幎y/����G�|˖�~��T�lh�b|2|��>q�=Y�w��Q�|����dM>FV�I��L��լ.�� ��å�>&�/Y�����aB�2��4��E8
�ھ�ԯhy�x�$醴%,���Qur�QfZx�O=N<�P����;\�璧
dL�W�gMw�̎�eR:x��e�0��_=�fȧ#V؎χ#���0���G�O��ά�F:%+#�V��o9���"���}�k�Q������ط}ÄH����1��tI��V�m�ǅ.���(��@���h�ч��^�!��,��y1{-�\�}/��W�1�v.N���yo"��^�z�i*�u�k�K�z������9F��s�����1M[Gg�|�T�L&�6|�݉�íjZ�ǪV�MZ�ܚ�ԕ�sS����z�,[����F��fNS�r<�������y�c�Z���>ܔ�*������˫El�IsZ<�2��l�S�y�5�gr��<ѬQ<uIk���m[;#�6s�u���+U5����]��n�GD�>�ݾ�*t���z�\ԾF�dM�7��|����5ڥ=8�=rٵ�1癞��^[U�_�]sw���R�3���^�r��沭ԗu��j��k�cϣ�s\�_<�����   �T  )  � �  3*� $ �׾�7��_��ף����yMUw*��t�*�^}S�\���Z�#2h[3Q�����:<�Uk��\���G����=q-���Ȓ}VNխ�H�:��W,k�y.S�����)��Zy�7���~GN�9��q�f�q��`L�%i}�Ob�Ώ�����o�k�F�<4�ɟa�cV�(���0������xj��a15ם��l�k�Q)l��L���[�z�ђc�w�^���'�Dl2�H�स�I�n��0jg�v�;d�GA���v���l-6|��wX.l�z�``J;5�!��GL�zQ��Ff�=gMV��`���>��s��k�$r�$�F�͞��S�����U�v������jX�����1�|;M<��`���ӍKϔž��e��k��k�����^�J���p�Τv.z0c���cg��y�K����R\�"���.y�6&u�|���[�s�u�x"'��h�; ���$�:p��B�}t�tf������e^��>ukq�?��\�M��=U�3�f�k�ab��2i&8x�f�Ν6tنb(��1^�"�Фx���c�/$:h��(�G���Q�t�Q��+L2ic�s\��b�yGZ"��b��:[VN�W?:�*����D��֛/f9�J�>�)�5���S;"��:�^�6UD��k%5H����n6;?Y�:�/qã���a��(���}�]�|²��.���uJ�Ee2R������n�!��<�RgjU(8}�n���dz��ݼ��oNS�y�ڬ�QݞE��P���%nH�H�ȯ:�"�tr�Y��Ǵ��|yt(pė1��]��Bg�<�Y�d��W�$�:C�琑Yd�!AR�N�F���L����P����헗�ذ�m�a��k:Ѫ��I����$Y���4a�%��&zY���Wtc7���g����C��%��o��:��x�Eɺ�Y�.dI'$���]��.�+�t�%ԒR��2���]�R*�S�B�T��V�Ԋj��usL��\�NMɥI����`���R�$�w�f�W�~ޝ�~��Ι�:gݭ��󽗳6gL��]����v�]��k���v�]��k���v�]��k���v�]읓�v�wd��rL����H�7�vN��;'d읓��V]=[p��۷ٽ;���[��h��7wGp�����!�BMDD�ɓ&L���fffs��>�֨ ����^s�zzwZ�  >�`  OL�2dɭ&�       �{�    330,�&M�����L��CP��f�f���q���A�?��9330���330jff�ff`,��,����e��q>���fffYe�X��������DM�DDH������>�D�ɓ&L����ٹ���Ȉ������������dɓ&DDDDDDDDD����DDDDDDDDDDDDDDDDH�  ��   �33  ;;>��       ~��h  ��Ye�=����f������330f�flg{�Z������2dɓ"""Y�&L��������陘���330fe����MMDD�ɓ&L���ٓ&L��'��,�w�Ks0���330ff`,��s���33fff�33�e��� � �|�hѸ�`~ ��޹�����vff`,���Y���e�Y,DDG���m�Y�����s��2ff`,���Y���,��7舙��pYe��&�"""}q��9�t�4��� �|�33陙��33,��92dɓ"rYe���@  zff`=330s���q���A�? 	��f`7 j�Nv����330ff`,�̖t铧��cQF6dɓ�N:`�-�����     ��D���   ]�m�      ���   ����5�      ��`    P�  �m         zfg���        �{� ,���,�},��DO�"bd��,�ɓ&L�̙2d�e�Y@    [m    �M4h�ӧ8&1�b�Y��������DM�DDH������������,���O���(� ���4�˅��It�/($�$�F�>0�7I���%��4Tx4'��0iZI�Kp$\!��D��I�ܟ}.��QUG�ьϑ\��b�,�a�#��$�VMJv)��ǲ��b���(��"�ɍn���K������H����U���ǯ-���I6�wf�)�ۗ]��a��7��S�.��^�=�w*H� �2�k�ݓ�zL�OT8*���l��sml�U����B�c�yY���W�1�]O4V���[�㕙��������Gm�yJKs�gnC�$��Z�*�s$�0��1_=�K�)�����nN�n�|��}&r[f�mj��]���M����Vs{�=�����|v<��su�3���f�<��V�]+6�^���Q��.��9��zs�o�o�b�u��i,+��zr�Iv���W���	"{��=���K^�EG$�էus�7w2����nv�Uͻ�ǽӭ�wgvN��;'n�܏ul�η�+��}����v��˻mݮU��uٷ��F=�u���Ε�+:U�V���j����]��Y�s�]��k���v�]��������{���ok���v�]��k���v�]��k���v��s������$jJ���%�Q�ޙ�������}Kz6���H���y�{��ܹ�wsU�6�<���ڪMQ�ݮ4���۩F��w.���mݥvy�j��m�>���I�����)i˭�FBz�]��q�Ͳ��D���+�i�����N�kq��-u�]u���7'd읕���f��Ͼ����vNη�d�w:[�rnR�m����.ٹ;'d���;gwS�Q��vnι�[9��*]%@�Y�I?�nA�'$_!�黸���y�ٗw�L���vu�{u�;HTn<�f�S�o[�7���M[���&Wj�۝������;�vN�ٯ^�����R>�.�&��Iݫ[�͒�c�띝��ww73w`�j��.V"��Vͪ�[H;�]O��y7�#�Z��^Ov���N����\oa�rt�����y����w&LX1�gc��.�C&j�����xu�gV:��Щ�%IP�u���Ů,�uŤV�S�Y��oz�8��r�qa�nսFu���k��t�����۽ݛ�;'d읓�iZ[k��ImM�뻾�%ƛD�Ȋ��ѡ�׶J�M67^�%pJ�X+��cve��B�:����<�h"�[EP[��{qmE�oy�2���;F��1�e[�����uֲ��ⱂ�E�I�u3���ظ�ݝ�S*�5���V[�F��WV�s��Sɭ�]�m��y��j�����n�+5&[ֺ�ǹ7'd��;gvK{o�Fl�K��G1�M�;'d-UW��.���m1��Z��,@͗�Cv�����[���ع�� �2���[U��m��e��,�7^�����r�U�s�3�t�{:�k�޺�w�=Y�fs��|��q�q\�Җ��.ٙ�tǼ�%x����t絻�{����U�U*^�\�����Ù��[ӊ�J_B������;��Ut��{������f���y��i�G!�ap}��\׊U��أ�x�mm�CB^!VHI��	RrbWw�dRuk=���)Nj��z�p�����Sk'6��u��grԪ��/���n������[}2�[K���M�с�4s�7u����:gBs���t��w�6]��;'d��|�7;_K��.��%��׈4��[v�Z�we㲠��W�*L;o^�ffk��n�-i$���;#�w��U(yUS�#x�'ff.��#%͓&��ś{�ٱ.F{p��V*��s;�ۤ�f'�R+�L�����R6����B�H�	��,��R��)%����=2g>�y7�tΕ�L�E{+U���f��Ц��z���ۙ����dr�U�&�>�9��v[L�\&gLU{;�
�wr={ӳ�i:���Ϋ�Y�^��:'6e�6�c��|{�L<j���U1r0�紇wC��x����3m�|��v�Ew���kz��b�w�G{5-��dz2S)��c��˺��۪�����;'d쎜ݤ�'��ޭ�3�tΙ3�m��Ԕ��ݭl�&2j���O7rvN��O��L�ɹ;)R�~o���P��N�K鏳w'd��)�ct۔��+f��wngm*'��t�m��3�;��{3f|�p���S�.}�7wf�Χq�˙�J6�n��������=Ź������9�z�������v���<�=�z6��M�1j��M��&�����Y�;�Vܮ���z�5���t��$I7fvN�}k��Ի{�j�m3��m�{չ�gk��7��w۶����omն�]��k���v�]�շ��v�]��Kv��x�[UrA1H�m���{���dݱ{�E�6�X���l݂I�ڻO;�nN�آ��$��gd샳��s��6f��?�$�웜�q�M�.�;��6�w"�_=��lQ�5�����Q�F��tSN��ӕ����Q��J���;hJO�{�fm�����3�װeDhoN!���:�S��<�gnZ�S9��"��۝��a�ĝ�vV{�x-�vJ���������ֵ^���0R�Љ�I���"�*$���9]s^HA�uE�V�ܼ����ʷo;u<̝z����lL����x��n�j^n����4�ݙ}{�3H#��F�`�]��>�P�n���Z����2��0��d��-о}�p�u�����L�[N�tVU�$"2��j ���������/v⽲����ԓ�v>9�wY��M9��$�Z��Vj��	?:J�%�"��Գv8�U+��n�]�;Z�q���MM\#Y���.��0H�=���_!�M���[�AK[�"��sl�m�0�

t�o�uY�Gs:.��Bv����[��'�������K;d��ͽ��0tޖ���-͝y���IWSOK.�P޽��L����!H�$4`aE�j��r��}:(]&cu��@��A��錖��H�s��ʅWO�N}ϋJB³)��bO��Q�fͲ�:CL�у9s%>�Wp(v���i��X[|v�.�k+~�6�̶*	ՙ��4��R��i��M�zU�L1�.�;�}Z�Ev �؎���j��~���z��[����*���c�%�d�Zq�'j36#���]�Y����BR�4�N�WX����9t6�t�{:�慯	�%	w�7���F���IWd�W�Bz�-��9o}�S3�f�z�J��;s�r9�/�F�Տ9��ӕ9�	F�<�=�Ù%�$;�;�R�GgWm�/%w���[IÝU�ڽ!76�B�gf�Wt*j���F�$s��n���7t���M����r�e���,��h�^�ڬ
KA���"e�물��]��vݤ^�u�Z��u)��2-%�yv7s6�[���]sۘ��Ȫ_X#����]ְ���s���4kW��3���7׍�h�YT�#��*��(���̓�o��1Pm�%�xv�7G��>���9Y�X�r\����Ŗ�֩�(n��
�3e�
t��r���.��ӛo!0��������;(F�\��-}ϲ�3�PkWUeA��
Z����r\2�c`�AC��s�EV�9��ڮ�B��5*�)٭	��<)���Ւ���ܜ��}6E�8���WכkfX�V�ZǤ��B����,�6),�b��U��K=\Q�}u��������n-bōk.+yeC��\tޡٗ�o[�0�|��ܬ���.�{n[Ӳ��9���Cr=�n�%�W����=.�*8.�n�L�w��{5�幽���U؇d&TPn�l�x��ޣo���m8�;M!�7�&�$����
�w���"�G6F;(5X1�w����C�^c-_{Al�ѩ��JPy3N��̉e�)Co�-��hȦa��k,=�X�侥9�nu֞1Y�F��o魩���M�6U�?Z�A��N�dZ�P�st弝���+��n-z�ؖ��sޏ�p�3Fz��ayjc�Ӽ��ۮur=���3�N��K����W/NweiD��q�3��s֛�i�6�~ޝ�em���1
�};z�7�V�V̨W)���R금u%���sc��������F<(��e��eSe��_*��׼OK�2vv4)�����R�d� s+81��鍆�[(VaC�"g��*7U nz�Jq9k�U��/o��JC2�Lpn�D�b�<�Ι�l����+m"xĽ�%;[b�l�<ْ�s��;�p$��)p�۽��:�	ƍ.s�n����
�3�ٜ��)*��#ʰ�[�߳�wwV7��L\��X�5gR��G��LPἼ���G���^F-��e�,Yp�������0e�7�U�|���y9OOS����R�w\��!ػR��E��VڛU[�����0*=���[��ط���G�ޥfU;j5�vt�2�%�B�!�é���O�RȺ���Xl��V��*cR�����-މ]m"��`�E������Sr�8n�6Y�o�%u��"T�U�հ�
sJ|+���e���{"	M珖�\wN�a�nv����ZS=�16su;�Mv���+��u"i8��r3V'�"�Z�
���k�'��șe���1�{"��.����r}�=N�6#��Ǵ#9�D�掬eؚ��d��̩�ٚ�7����gv����t��u�z�ݛiԨ-/v�T�{xYr�<��]JFU��6��v���%��Q*%%�b8��qD�PX��L��0��^�<tӈ�<-f�VA�ͫZ�!2v�}����f.�����0�d���Jt5;s%�nd�{2����J^D�	R��]�.�^=׍��؆�,�/ftԌ����yT亮�s&�e0˽�X��$����u��b���t�]Cm�:��.�8c��2���uxQ��3D.���.�ͱ}��_j�owܧ��vv��j�k���Zwz�k԰d�uZ��׻ZL�c�f�e�Un�x59iS�8jK���oz.k�_h��OغB���W����޻gx'&��{i�,�D�w���:֯�lUo.�;�[�y��֪[�ݶt�b�l��9YjRV���Cw��k
�I�k!�JaٹC��:]��8�D�G�:�\��j}l����=˻�An^o�*C��=u�N'�#s�Ww'Gè�	|�q�;�)���;�cv>�q>��s2�"����7y�r����\�z��wA�������+r��ʌ�(1�t�vf>5��f_�`�:�zƻ4�ďj�]J�Oi们�Y:�\�,��4�$�C)W�,�,��2��0q��C+�J:K'm�5���R�ԣ��Op;R�sx�����'9uc�Шt�Ν�_\op���7���ޠ�ɵ��4���N3�]1���Ψ�3�`ꋷ����J5�����x�w7,���o:��d���b���f<��Z{Kq�z&͛}V������akʷ���Fm�7��cv�m]Wl#�����K&�n��-��;.I-vh��D�TV����G�E愤4"G-�����Z-��:��UNT9=�{�_��]dH����Dw+5u�Ցm���Ey����ŷw�p��͜�wԾp�'�g<q��?f����T��MC�M�����v��k|�qg(w��L]:##�ݛ�n6�=��>�B�S-7|]��©VN���[w�ǯ���|���Vj�0X���]��,����QIQ�#(̆T�F�	����.�pN�(d'/fD�B����j��bqw�Ի��޹F�p���or�6��]+��"�R��`��5��^�cp�料U�]m���Ӧ�8�%ٝ)QҶJ��9TSf6C�j�4����6ދ��ֈ���;�S�ަ�F��w�b����kg��j�Op���r���A�C�=��7��.��)͝�]�e8#p��c���I$��c����!$ ���� C��	�����~������p�R���&��3��O��?��W�~�������k�/��뎷��Fv5\5Ƴf�g	��=t�I����C�$K� �QbJ�b]NMV�ӂ�6�i���&�<�(�S�-�ս�hOh��c=on�
ڭ�#�D���G$l~�K������ݩ�m=�k�dى�F���Nc������J���7z��H�U�wH�Q������M��{�aPfW=z�0cR	���^m��۝]X^�o�"�>��7e�����������_WD)��{m�93c�3�[n/f�g��-�:��;�K�$��!V�Ǻ�BV�};�ʭ��/7l�����Y��xA��L���twd�[����GCs��!f7�LWR�U]�N�E�e�����d�"��I a���eJ5���z%�C�q�x��sq��ӕ|B��pkV���۱+C�S�p�XJ�2�9�t��@��{�۩d��s:��Oz�5Y%� :ܬ��H]�0umq^���\�M0F�P������PM���]�mΑ�P��f��c�����ѻz��7�!ո����Gqu-��sp5K{x�9�[]�ٕ����"V�o!�4�� y�]����
��]��9IhtNFe��q�T4Sk6m#z��9V���8�(�En��{\ho�����gM��nm����������rc7 m	��k���F�M��4颜�#v5�U��+z��\:���A��2��R���b+��MԷQaC��Rn�I��]�{[Ӕ�t��m�s�jwl�l<�6���W����I:�7)���N��E[[�����^�u��3tJ�!N}�V�ع����n���ވ<�h/w����.�|R=��#���yױa�t+����ζt5XTT������\�f�BȾ7��U����={1�49�����3��T��c���Dx{�7L�tv'!�n�:�ܢ�E[gƍ)^�6��'��w��-p����,�����靘�����Q��h�c�_R���I�`y����]�F����i`�ImޱGZ�����k�m�U[��r�Ȏ��}��tO��4:��u��t;�;|�L�j���ھ����H�A�}�V��哖k!��T`�mn)�����e���Y���x6m{[Y���R���N���Z�mrR��Ȑ���W	�M������̝x��t>|[�KW�!�O���)��| X�Ǉ9��̭�z�x8:���),�O�#o����s|�G3�2��cY8�ʧ��[׺��od#���Jӛ�z���6�{�Q�)��vѐ\y-�B��2���u9�:�n�v%��v�� r���}��N���Mΰ���,J[��xa���b>4yc�':n���$�̏\��6gs�.4)��RGP��u�mܝVg]�c���o&��f�]t��SC�ɦb��� {��� �T2묕��Λ��Ӯ��֥�+˗4�y�gr�ZssmUo<x�\���H钬�ڔ�m �1HH�
���o�!3�����%]��Ž�⛦o�)}�㣃1��L��rQ]�B.�r)+�<�ۭ쾦��v�����cN	���olG ��H�H�r�$��I4j�Y�oy�����p�En\�s�Xt�����n�n�EK��1�V��j��z�-d�ú�GoN��[usk|p=;iz�]gS�ژ:�ڡ����$�U����뵶3S��(e󋮥s|B�r6ʱ	�.�<x�twe�����q��̛�W�r�F����[����.����+��
�s��rT�z�X�[�KjnT���4������5l9�b��c�N�.�pm'b��X���Nڜ��\s-��%�a�A�z��C��"����{cf�|!Y�7����f]��{� *�U�����v�B��[wV�r�ӝ[�����Y��hѤ.��Xh���{E��<:�%I�&�������2��[V����%ڛϴut�Liռ�.�_	-v�P��M4r��,v�nɹ�\[�͗�]��3�tS��)���5h��N5aPg}t��՛G�F�C�yz�֯m��(��7��{�M�ʸ���oW�V_tA�c#>�]f9��yz�`��`r�KP���h��e+l/�N	�J���W]���@�rm(�dYN���5|�Z[��Afnc�ޣj�M����G�Q�[G��W�ۦs=I�E��Cm^l�}���4]��G�.��+4 m�q�:�{�Z9ݫvD��.�1�U͵��Y��١j��ޜ��xۋ;}w��c�$���鄚�3�U)�n�j���������5]�QZ��Z3�Ҹ+%j���m�e�Ѻ�Ó�2��+�Z�F�'�o���O����ʦlp)�}�N�T�;j��3tq3�J|j�	�ޏ�]4D�1UX]�,M�x-��wKd�<H+Er�<l�CTK���v2�y����:VS���y���g$�/�G�:���U���б��b��"���Z�}��w݈vd�]��Y��ml�9���u�6��A��z��S���x����m��յf�f�N;�{2r�4��m�K'v��WjX�յS]�0E:��������:)M�Z����S0$�y�U{�* k�w����ݙp�$dY�ء㪷�L�{/�A��|<�+�%s�3F,�F�sM��h� �����v����wx�ʚ�����g\h�!+�b E�;�����4���:�t*�ӡƟ=�4��.�K��[����|�Ǽ�;Ԗ<� Y!���kZƓf:�Z�g�f�9�{<Һ��Ŵ2���m������W����C�v´��9I�Mͼ݆=� <U�ȓ�ۙ�YM���z>x�a�[���B�!�vf1,@�4Ք��- ��$�a1�l�$� �;N���:����4��.ޝQ߇�e�������GݤrAǌٽ0�����kT���kWl����&�	�oN�T�%i�lm�aX�BS��>CE���Ǥ=�W��|t��>B���8U�3;qm]��ٜU�a�U���jp��7v�1�燷s)xg�0�j���2��b��E��۽g��k�SM�s8�Wj��鈵�uVI��1��lᬧ���n��mo>�7������Ѵ�v��R���Mk�7h�Ye-�yΰ����.��3u�!��X�	g�a�R�ݸ��Cv�sT�$��SټDt�|�׺��D�m���`�h��w9�5�C�a�l,�j�Vs.��;{�lB��7t6=�5�P��ee��S�C,@�\(U�tq�N���J��V�o9�6p��Z���[�XF5����L�|���n����kxjh��Zj��<y=9��^����=�x_5t.L��v�UoUV�\���x�_auwj��9�M�wt|�!���ܹ�K��Om���}Wn��	�y!Bݥ|�w��z)���CI�s����s5Tc+j/1�X�/ ���̞E����NT��Ga\b�N"+ԃ��Ɲ���ISP��b4�f����Qݼ�|���!(��3Ov�n
�XX�n��Ka��YG�ܼ�T��e��S�;�մV$����F.���WSJZ}�b�KʩKN�8��C/�\��\�-���hX��L�Ś!�1���Z*�r�5]�e=d��]��n=�myV���]��nU;_^ǝ{�	u�����t�gl�vrS=�����'« �b���/���BG��"��5uH�p��R3U�7��r=��@��,�z��z_K��_b\�t H��U\P�z�j2�2�ᗛGyt׷n�h�����O��՜�TuϨ�Ù;q���hUK��=9c��«5́�qmʺ!n��z�s��+���OV��mQ��7�K��OK��m9�A�ƽT�,�ݾ�Ǘ��UU�{��*9�g��f!�,��tv��Ұ��Y�s �����	v]�DzHz�Rqs����N�lX�����ԁ���Gl�E�X*� s����!%.)�\*TƐ\�u��mN`C���x�*v�@���dcJ�Vn�{� ����N�X�n��x�D%�B�W<�]
���.M��.˹���o�u-F�3�t���6,�.U�Y�b�s�ˮ]kBwc�������*ۣg[��
6-�2�]-�Ot�§[�j�auUJrOB�]��kx�xx
�j�Y|F�=s��)�>��V�M��]:Wr��vڌ_,u��%r:��Mpq'�������+��[w��@���
����6An�:�kr<������Z�ݘ��;��  ��g���r�����$ �!��z��q�B �B"@"��8�q�B�"� � �H�F""DA0�!ȄG�s�     �B9�   �     ���                            9��"$���A��#"$DPFD!��@BA!�p�B �D q��!�Dp�È@BA@�#PU�
#T�RU��� �"�)�	�����?�n���{�߀����������������T���o�־�f�ss������9�Y�e����Od��pӽ��ODm�7�� 9{k��D#;y��>�8�(5���]��IP�נi$��&�m�~$�P,�6 m�$�!2@^�@�[�m�KmN�d�6�i���ms&���ZD�V*�����$�&��]4���]��[���\��r,�'zs(S�V5�8I�;��l��<��\z�x��"�b�nI�ݗ�`ЙrF�<���R��
]G9,��7y��H;0Xè`��gj/e+��t2xq�kKF�_X9�N�wХ!2���0`�yo	];R�����+0r�YD΃��١=��Z��V�9��+���u"�*͛�-٤��D�$��;/��ҳ�,�u"%Q��ѾH`�Y����.����w���,��;�`*�W�}v������&��i��F��/GU{n�ɥn'���Iwiۮ齽4'�o�|��{z+窣��'egtպ��KI�5�I��v�m�*��y�+U�k^�[�X��w�V���0�9�%�7�e�,]%y�j�f���r_t�$MKL�D��̦��!��<\&3&���^w.S/��g7+�=��[|��NH�*C�+B�|~��9�A�6'��9,�XAα ,ɾ��$m""���'[#W���,3N�#�o�;�TF�'F�1B�r�݂ռo_?&K�$2m�*',cZ��6� �V�KVu� T���Q	$�VV1X2b��%r����q��{�3E�A�}=���y��dU���e�T��C~��M���yq>�f*����u9F�2HŬ,J��T���X�6��;��G��+-6���#�b��UK7UNb�[�
��cc�)��ٺi�_�*
����R%�M��+��[$��IZ��ў��ٴ��&��!Őu�N�klĽE��Pt9�L����LՊA��t7�i�p�l�R�,�T��_A��ڬͣ��`D�J�E�f��-獤�����tN�p�Q�+����9(�������|t7hv�8�#�� ��L�s�>�7|���]���Z��NHÊ)m���"ɧ�MWO՚p6��wb�c#)C�������Vփ�m�"���[��g93�V��ԃʁL��A�ԭT�Z���X)�p�1�oo��I&�A��_�8�����ׂ o{r�3�͝>��Z�'n:K�*$���/��;�+6~� pR���)�g<��:�^+�0e��k#�g�u�,���؍dA�	��ྏ
��E�e�֌ PxJ�!�"���c4͑��5�N�ig�;���4F��Z��=��^��B{w�5���wHګ�%+ 2��!�}�x�^�d�d�/9�4������\���wA	�D2����l�0�PO�����5��t/MA�9�ܝ#����>a�ى$x�!G͔AY�v��v2�>�'�����A� e�	K��s���_�[��£�0����;4+�����}����Hg?����=��}���C��$1k��rvv�%܃ht�P�Ni���:=���)�
�0\�Hʩ
T��)��a˫��uS-oz/y��\�" �#���N���/�@.�G�U��]L�;�e�a%�>	�ۜ7�7\�]W��|'ܢ�YZ����qW���m}M��/i�h4!$2�}�h6t�����ϫ'|�m�B�Ϣ��� �W��+�x|����kM��I��:�_[H�#r�}H�^!�fm ~���A�NLr�}���v%�󷗶��U.�K5HQ�������W�����#�{W�2�p�@{�����:��0P�Dw/:H�Q�C�!=Sn?��ʆR�`ߵA�8j��zLX@e��>ۦ3Z����FZWRl���Q�X}�Sbz>T���m�ۼH@��W
M�|~O���G�ۡr�n�y�]f���U��^���35F켮qv��ku�`�4SBU1Ji%�(B���)"&X"�S�^���H��݃	�B1��|OK�@q�<wu7�{Z����>�N.���>�8�b���C�*#�
A�e(}T:NtϾ�c�ٻ��I��~��覭���c��9Nꢛ���Ts�k3�'3
�}w�IYU���NmH�Y���'���/�N��ז]|"ߚ �̀�KE�k��^���}]7P-%�	!���O��ىB�q�=�j�X*�ۄW�=K�Y�R)�H�>��e���o�u��{��j׃����Jq3�x*�\ot���;$*�I%��(�������x�}���{���9�Z����[37%;�:
�dj5�ȢkL���n�K�4@�F�%O�����0`|�Q�ڞ!$Ӊ��!.8�M��m3�a(X��\�:�SHSf&�����Qe�0��a��n�b7��8/oD��L�K(�NMO$���T�=����w�ܡ��zZ���H���'�]�M��m�����y�}&���z���E*c	՜��ҝ�i�������\��5}t
܄���_"s��=��?xz�ZtN���	�B-0�\�.���c���1�{}����ݵ�]NʵW��J��G��׽��죄�
�0�1�C��sV}Et���xh��z���վV~4F��>ؼvTy��|<+^��a��O�*����O�K�p���i��{�xk�L �ܛd�Ô��꠨���}�"�i����e�ar/��Hz;�)mY�V���i�FlGf���_nw���(^.ɢw{~���8�����7P��֯~E���ER�z�*O�������w�hV�ʾKD"����R�Nn(T$>f퍡anr���y���%����Y�������4D��|�����GkB̺)���z+E�.�ϫ��@���4\4e�AYh�v�[6�ĸ��*h�ou��Uc8��e5�� ͯ�;~�g��#�/�.�◽7�5����[՟O��P�w$�)���*�'�zNo^�t�NW�`�3�5RYf�U����脏������~��3��Ś�`!��S�������Hl�{�����N���	�s]�,c��:g���5o�n�_.2�Ld�'���-������ea8�N'	���ޱ̧�bt�N�f!�͟$p�D���eX'秾{3	z<sE��L��t��Q],>�Y����gl�z//�8GZ�n�1�-��}�ͫ���8�O�`��g��b�Խuٛ���
�؋jg���>#�lzV��gǫ�n���#a+zr�WӸ�<��E�gl��Q1UdR����c��n��n�,R:�GIE�HI nr��}
#�J��AY�I���t��/����no|, -9�ɜ�z�cns]n�rVV��� Ba1�u�M��B�j{��'���P�f8w�L�rcm$������
��&�DtK�*8�| �铭��Aۦ��kx�I~�]ա�ė���5��I����T��{�I'HQ�ߒ0�� t!�n|<��!��L�oke�@�!���t1�;W���(��χj�F H�J�'u��e`�u�][M�
��;nm���({ +8Ed�`��m��q�5�{7x߷�� �Y$��2�L�Prz�_���ύ������b��r����ˣ�G��
�Z�#���ݘE�^ϳOt���By:�:9Y���j�/,�!2�V��[���kҧT��z	��dR��H2��p�E�ZZ�U2g(C��	�P�,p�|<1)?~�'�}N&	��<ϲDM�;�a��5�o]�����S=�S9�5�޲f݄Y�޻�J|</H�Z1#A"�Fg���^�W�
�u�0�~�c�H+���o	���ͻ�{�>���!�d=���hGG��S[�j�͡vq��a
��r�?q�����������Vh�D�o�u�y]�'k��p0��oԧ��z�Eu�*��%���q�g����y��p��x���ps�uuRB>�G)v��	�dʭ���Z"���C�s�}����V�۵[��G���>����pQ�h���/�o%�7lF���*���ٔ�[���w\0`����q��Zq�r6S)2�۪7l�����08Q��CTRH�q��_"����*�{�6@��/Y�x��7^��j��aKY�Q*�KTp��Z!=%cLu]��v���#��mwn��j��I)$Ea�����v4�Ś>�Be�>ʱPt��rR휃{���a�W�����}\� s9:Gى��|<$�kF�ŝ�8��䎓t+�>cP��t�������I��}�9�"�
>w��f�C}�bd��j�,@��;	�x���U#�>�a��y]�	!��>8��Y]
��lc�*�6q٭�}�McE�i��&���=JM�� ����)�l�vm�!E�'�9�R| 6A���Zf�1�T���>�+z�,�#z��Hկ�.�>� y�?tdqX��m�o�M�=w�ϴ�'16��j����X��|#'�U(<5ܚ�i�|Mi]��7{�c��X4ha(�V󫋑RF��De�kzݤA��CP4�!Y˼�����	c(�FCW2���n��X8uv��*ǫtZ���h1
�y<���x���&V'-��+�9]��Kd��R}���U�?�u^�#���Zf�2�f2M_/� {�f���|^�WD>�Z5E��T=�U�����W>{��1MLZ6����U2�|p�}�Y�яS��y�z׳O�o�0�Ӗc%q��C��Y�xz�S~[��}�T,��f�5/v'I��bx�9�e��
�����z٭�[3��쮐����j�:!czI��}�b*���@��>t=� ��_�.dX�_}�=������1�kYsYe���0��	�svug�3��,t)����,;/!\��K�o|�(d0��x�T�ƱZɌ��
�`�)���Q�����`��1J�I,ա��i(D%���+1�<�(v�T���u�n�ʃ3S�7u1��Sh�Q6ܛC3#��L��d���mY2y6d��z�k����������D��:��J�x,v��^�>��@��+T��h��s��u"�/=įt��O��)���wO��Lgʱ >!S��8�e��T�M�q�}��Ԩ��J5U�n1!��U�ƈ���{�#��� 0��Эz��d�1z����e0!�PO����n��g�HY�k���2��Ī��ӄC�r�>�c���86}��U�4���"��p_/��G{�[���`�eZ���!R�>��F�����#��1�4P���!w�L�!c䇔Q��~kOl�k*����f�M7���,�E�F��h�@����>�_/H%�bt2vP���q�ȏa��.�������t4�0���a�H/�#)8p��{@@�|����@�X��S{y���{ê��t��toV�oS�I�%�{ڶ`��R�+��K��a�����|D��nǒ��M�c��C�R��'d�Hg����2�=ټY�eu�	$�-p��w*)3&`l鴰�T���=n��̩����BQ�gu����yv��2��^����U�R6� �u혝��Ev���͐+q�+��Sy���U̘��-�lH=�T���������ĭ�[��Wf\=���^�M;��KkuR̨�J��v�|Wf�i]z�ֻ����o�}���>�
;���lyK5�ȩ��v.�RΣ^��a���a�`Gj���fk>p�˝V�Jm4�!�BWr���n�u��6M2iS)'�i�e��@0����ƌ��(q�(Go��}�s���(�.4I��I���(�*75������|�w������ ������DD���DDDDD~ ��秥������vvvd�-��[A���n}95>�65 �} |	��}��}m {�� ������gf�,�&DD �
��v�J�@����%��B��I6�>@�a �daĈ1� ��	�%��2H�QDLQEn���&"AB�� �L��R�&CA$��������D�H��$�-쐞Yii�(���Ϊ{Y�D[��R*5��0V��P$�D��N�c�8�>�Q@�
8a)�Kt��Uo�ʇѢ��6�ه�a6"�M��TZ�4ъ@�&}��љ�Ճa���0��
�2""I�����U�U���j��)��EwJ5D�Q�l&���w�~}:�����Fд���=Sqi�<��ڛZ��D��ݛ�͎��w����Z���\6�zà�fl9G4\�uI^���X�Uy/i���<:[N��U�t�{���"	���4����'�rj�]��:��xE�Yo��->�<[SN�[n���G�xgAǘ����csR����I����z�`@�IxF����ю�m��=�4���u��Ԇ�G����*�+�[�e���Z���R"�-�u�n�zXxd!�W�v���v�,�%��vm`a�����6���H�����ehs|e�3����#8��Wgo��y��SE&��)1���@�0�z���B�^�ˬ'�j��l~�""�qsWC�K�Y��!R��d=�X@��yZ�{�ʇ��Zىɷ�n�D��B:#��Ҷ]�o9t�o��E��%]^���-��,� rLwbQ;��\�~�����j>��#*�!n㷲'^v鳖P6�.9ijQmna��e{U��]t�S[EN�IP���!��U�'��i���H�ݕ;(�5�ں�)�չ�i�v��wK����4܉�h�gpX):���9�=;��Ca8nU�@+o�b�4uQ�gOg#��E���!�%�%3�cGq�f�&��M��+CZ���vZ;AH.)��c<ڗU�H+���X�0�L��6	+[�y{i�����5��Uݖ����%�<��PF}0ǛX���=�;T�R[d�B�p��&�nz��Q��޺��_����])r�:�f��|��ݵfV��c��Z�v]v���E!Ǥ5�������1�d�o����
CL��,�jH�j��JCIH,:ɶKAH
j�V���M0ۇ.���OR
C�%xkm{��7�!�q&�j�2�R��0 ]Pv��U)��)�R̜Bؤ3T��%k;���������|�Q� u)�	\���i��@8�����Q�q�a �(�	�Q5��d�E��9G4Q���s���c����Ϡ����
C	1���i��m ��R��h,�C̛C��;TAI)����=��VZA��#���xQ ��i��GƔ:�_L�PR!)r���lb�i4��m��a)4�J`(N!�|s��{߽��[���TI�	h(,$Uf�-���u�[����3�g�d��RAE�e��<j����*���3��}��~{!�@)ݹv��0̡���CHZ
CH�R*�l�uP�KC,��H�)�9�k�h�(��b����̖é�k9ɴ�RI����

a��C�i���`-$�'{D�b��T�6���Cy5�7�� e��m)'B�P��!�5L��)���M�*�I7��{Z�ؠe����6�C�E3)%����~������u2�b��'���C6r䤊!��Xb�j��2u��Y��S6�$�@ � v:�K�J�n���N���n5�L��Ac�i�Vѻ���e��1'AE�r�B+�s�ٔ�ݡ���p��(-oRL�����n(���P�1���E�A��H��������q&HLd���1Rw���v��f���uJ�V3o96U"�6�� r0�R��Ϊ� @��t}�|5�@&�R�̴�C�A�)�X���Y9�@q�"�(r�T8�`[6��b�0�C�N7 �I�vU*z����Y��HB��R}t) $�ۖa��I�h@�hP�`:ɞd���*�Zyx}��w^�ʳ�AL�-2��&�8��5V���JAa��Rp̡�ي�.�-!�-!�
AgУ����^��d�(T>d>L �m����Ī����4��VcyR�OR
C�@((kN��ha4��^y[����m��ABm% ���W
�	I��2y����P
C��0�{z��� |Cz׵��9��e���PZ
C,�����Hi6�j���l�P�ABkTMb���Kc�Hb�����o�o�z!H1$�
XRiުҙ�II�R��h)f�hy�gj�()
AL��p��I4���8��h�=_b�I	5���l
Cڻ�gT[��[&�_*R�)4�)�C����H]Pe&�-�m�1�/��vH�|� f�T4��}���
t$-�@QF!�O0�Y�n�JH
0��{�vn�g�fbA���X��ٽ7���A�0�CuA������) b��J.��e0���% �c4B�b9����L0�iMv����n��mi�ޮR�oe���m�%{N�gm��C��4���/ ,f�Fo�)$�r�'�����`��z�H�����!�5������B>�Q%4)G0k�ߝ�H�>W/���<1��:���X�I����o2gO�C$���$�h���H��b�i��ˮ���y)$���2���<�Cy9������h� �cTB�cu��4���'К�^�٧�-�1��!��yb�� `�$޾���ClR�UcUx�C	�;TRi$��R@U��k�������7�9�U�ۅ ((HoՆ)&��A�RP�kڲ���$�E ()=fL��CUA�>���Nn��|���� )�.�~��)"����C��6�R��0�C�ɫ
J}����)>�u�<�@K����e�(v�2����JR0�`�Z���oxވm9� ��%�{ǽk��>1��qF�ZT�'R
M!)!�Pe��j���B�R@���~��KI�L��_=�w��!��������"��4�ޮʾ���@X�7T��sD��m&��Pi$�b����7���J�*ڬc�s�?Y�8 ��JG�
J`.R�:�Ĵ�j�Pb@�M>�ZUQw@���6{!���g9��Q)j.�fh�D}��$/�C��
��b
Z�i�iHa% (9�@��!Ԙ�B�&��D[x���8{ȇ! �^�)f��q�g��()
AL��L e����E��)$׌X

�x"K�v)���{��)�5^\�v��v�ݹ�e^vt�_8�tI��,
0���?��>%�jK+3{�.+�����B��z��K9{E,s���:��Ʉu�Xw�,�y�3�o�)F�׉����qs��W��w&||Ah��]Ք��i
AM0
b�ߨ4��(�TI�AAd����К-��|w���JCw�g ��[{�Y�H
(�0��ݗ����@X�q!H7�!��a&P�Pe!�1͚�/�w�o��
C� �JLrQhZJ@�zQF3`��J׵��/�4Q� ���z�����N����>kw?1,�z,�v�{�$��r,�Q���aYj�i�Ƭ&,5��wn7[üe���S�,�'T?�f�9�!�/���*ފ��{�2�Ӎ4b���|K�Ӥ�I��w�t���6�Sg,����I�H[����k����|>b�^"Z;U��б���)z\;�I0;�K�6��:�	A ݗa�"�!��a�
HCi���4m�i�A�����c;���D�Lg�oӍ(��g��oL�e,���֦�yҎm{���)$�cfh����j�QH��5FM͊>��Kt�!Ń[B�:AE���q���Zp]��-9��v��q7�^���|�l{X�����v���A�WJB�MYIV4XؔR�.�N���g�h׬�5Y�{zI�LWu�$	dЩ�.����\��X_?1��� c?!;Ǻ����n����5n4�ȳ
A��<z��N��Wi�K �7 ;���RT���f3#��ͯ�/��l @ܻ٪q�w(f3fq�+7RϤ�>�J���o\�S�x��:�L��\�x�%�����9kz��U7�-!�<7�,�
�j��"D���̝���ܦ޼�������%��IBe�,lbU#������a�1�yϫf�&����Ƌ�C�<ɫ���0Y�ƹ�c�������/4TDC�ɕΊb��V7>c��t��?x{D<����U�����qI0)`�S�bE���K5�oZ�ќ��R�y��W��`���PϏ+x ��B}�{+�Y�K�,8��p�Q�"Zflp����B"q��l��H"܅Ga�)ֻ����vYMI�tuLTf&�l�a	���P۩�hӥ���W��ݱ��R(.O���"�� I��A'� �@6�����9?�x�Z5_X��b	�t��O��bZ���R�(���u����lEI�(�L�}{���{vX�3�0wZ��3d���n,�;��
Ȁ�G/D8��&$/��2�+�����te��3���W���ڒL
`����ِ�F�L�_�~c��g��HΚ�нH� ���T��	��1[^{پѽ�8�wG�6����y��ꂭ��4�`0��1B�v�vO��fzS���C1�3���Y��{3Eh���7��7�t����	`�:����f&[�5R�V=*�W�4m�y�7�>�Q��3P̓5˷���@�^����P��? /�;qآḱ�hg-���Ր��8Yp�4kVX�̶V}��`����s�s�+ѧ7!(����g���n�Ni��tޅ<�ͻ5�S��҈���|���e8�xx��H�+;�g�j���u�c:6�hЖ�E�le:*8[�%S����8��WiSE2R)#S3T�մ��W#1���{2
�7uʯ�!D���lT�ݻ�j�E
/����ɣ��PwI�@ �|sm�]!���̸�x�>�k�xP>"G���-��)x6'd���֘H��>�� ��2�B�	�5�Z���m��p�[$�` ZCI�J!��oA�ز�-��^!�z���9��]�с��غ�o������w>���QR�Y�����N�>_l�ݛ>���oo�+IGwe�9�^����%pH� ����^�1���י:�Q1R����
2��Yfj��ǳ{�3�-�-#X!�t2D� �sQftM	�\�Z�)�>�㩓et�wiQ�"����`�HL���r���x�eta�ːD��2hP��oU�;���eq�lĳ�s�3��Yz״�.�Y@�W=�z�:oo�^�m�7�>xag'm��k��t3DR�FESlU�Ø�w9��(}������Ӌy��vnja��Z��Nז��UF$ޭ�X��΁�	?�#m�������i��bd��6��%�+�W�&��k�j����{{I���D�� �G���#M��|�@������ubۗ�j}��6@&IXe�a^B)�JD!�Aˮjgތ�\=#�D�Ay;6n=A�����=+��cjOI�Ɇ�}e�'��y���`��7��@ن�j�b�p�ɥ6{yw����=R�V]���Vw�,�B��}�S���:���w$	��f��Ɗ�1^�F2�f�jԖp�Hc`�#o�፻Z3��j�s8��俸����G\z��݉�0��e�[-yYp�Q��?�����Qc\�uݓ��OxA8.�6B�k�|:7E����lƩ�����OdL�}d����.�[GS0ڐf�xc@�)y��ͧ�?{�v��(��E��sh��Y��w^����������D̉Y�*lƋ�����	�tY�� ]��zTqa��_=ƒ�
4��?J���;n�>z�:��	n��_WHH�����&��ŵ��ʮʼ�ؗ7�L�z
QV'`����i�C�<�ׄ��M̑o&EeQ�5EF)�JF�iz�0����a�Q�3y�"P̜��&��-^;�XQ��a�o������+/0}&�:5ƫ��ϨװgY.���F��rg�(��`���{ց�S`��N1^���Z40L��z��9GМ�z(�n���8iB�>�W���>�g�X���=y'
C|�� j���J@���ղ�W6�h D@}������C�x,�8B
�8nF��0` ��vk� �b���=P@�	�������o���3���Q���u�^��^��eDD9�̙Ӎ��s�/�s��%p��.������ ��$�2)��w�^R`&��LH�Z��6�*�9�E�ӆ�	�������))���6�J*E0C�ӎv�.�Tk�khgeY�Y���ϖ���MZ����_ڡ����%�boX'������}���K������?_%���U�۾,X$>��!N$K*Gm0�N8d�� 5�s�dIl$�j58��"�Q�	����)=�����ٕ1)�7NK��H�C��ϕ���L�JIK��fa��"�%�9i8ͬͿ��>�<k�X�3y��Z�{���9S9�w�.̰�G�=��kW��GJ���&9����n`�-��f�G>׳�tn�(C{ވ���(+w~ʪؖ���F��q�]0&�r�kX��T�,��>�3Ծ�s]�{�0�����v8���eɑ�0��ۈ��a�|<�u7`f��� ~.�g����Eѫ(C�ֽ5N4n��l��9����8x~	2�vW��O�f�e�>Ǎ}���A���w�1#���;Q����'�$�e(ܢ�f���l�5��c7E@�X����}��>!#$�	!��7��_��͜�G�(�[��(�F�e�}G�:�V�Z�6d�2h��Q�{��;6��\�w˝���T��5p�@�y����E��p�ó�_|5x6&4��A}�̙ӝ.i�Ie���8S�^�����n��V��4
�ڵ��^K\U�M����a�2*����s��Y�Gs3tԀX#�j�����x���/|�A���N�Eb�$�(CH�a��iC
h.�&q�`e2�i�'j������鹺�Ԉ�-�K�L�)`U�Js{�
!iP��6�L�qU���3\����ęޛB#Z�^�d6��k���Z!
8|1k
�n����hH��W�2����2;DY�[��<�������v��,D�]:��UG�Zi&l����^\\��$���s�S��ըMC>}�$Z���4�-�f�C�0��F�*�vu1��h�j+u�"&��xA���hT���67u�c���·RV=�\m��^�����x��N�r����C��z�����൯,��i��'�J�墐�;]��2ض���;Sg7�զ�������h�wW.N���\�uVE����-52�S|<'8&�4�1<qB��]�wq�����w��E�Z��Zȱ�e2[D��p�s\.[�cU�i8�P�6QJi$�u����C��N[;��������*c<�Q�0��0Z,���� ���u�Xߦ��֕�[���)g�V[<HƊ��ϴ�,�*ޤ�.��O5�]q���9��0�e�$0�	���%��r�o~����F��6��NOOK'����{ &[k���M}�5�s��33�Ye���=�z�;;�A�[C�鹽f ��� ����I���p%K0򋸾��g�UP�$�E�CA��D��R	��X�9$�R��d��.��*@ӄ�����L&Ӊ8"J	(n�bv6�����%��ҽ�T�6�F�p���F�o&�����f����`� շŞ�Z/�=��;��ܝ��g��Q�Zk�m�!4�A`��|nU;Hě.B�����IwUT踗ehZ���m��	�fbv�ⰻ���C:g
Q|�t`�@��6c!�oJެ��,���#%3���V�wm��B���/nUΉw��G^�;�e-\�W ]D��ۊ��t����+-�Z6�0�	Cp��Z�-�z�=��ɗ��Ens(�XgT��əD�̴�u	q�[T��y�<��%=��(���wm���c���K�W
µ,�q�ۛ2�X�m)/{�v�f�$�V޶�)���/�Շ݉�ݵH�L�K	֯6¥���3�y�6]z�e�.{!,m���+.Ne.�v���ˬkכ����7yD���aػ��p��<���R��NF�QF�Ұ�oj7x��;�J�6/7���}6�^���]+t��S��qI�
Z0�������Oi�>y�F6�_OY�5\�y:�ǹvqH�V�5�n'O	�Q'E�,W%��{��٨�ڌ�m'���]N�[��:�!�%]x1�5D'�
� �ܐ�̎�B"�=��i=K�H5&\���%N��nA��+[T^5w��8��yr���g�qOm���2�Vew��lJ]|٥���v��K�(nƂ �uי�T���at�`��X�qX/M���A�R�D�S۷�fx���<P!f�^	LP��A����w�Xu	V!�����Y��θ�#�_]1ĥ���p)�\����|��F֨�a��v�^�e���Ӕb�r�齰QZ�Vv�Sb�U�� ����f�v<5��M�[cu�w.�n�u�X7my�,\5��*���y.Ab�`�8lÐ�N	(�:�A2
�T��[$x  x(&��w��\4!�D+7���Ԍ��n2#�{�X�M�Vv��J��@��m����UY&�b�ۛ�L^�{�Ke ��p�Z�AȤT��[{5�X� ���T�i�~A6<�ȠI<kXrY,�7�s�C�똞���Z\
n�Y�(=G2is꬛��V5V�D3��^2?��9���� AdyG2	��z\;��D�[Y�ؿ�G �i���L���8�Iu0a������=r탄T���E/D8��&$/��2��
{�S�O��+�YC�`���.f5#�!mt:D��E�E��4��p]�����
�p��z.��{��jB�xS�wtt��N�E���s�3�h�*&�3����n�W@&��0�h_�$���d��v�$��l�tv�絮�S���%1Pv��N�����Hd��Q\��e��}��:��LyE��3�Օ�������_ۮ�=�}�/)\�V3`���e�4�('A{2z0��z�v���u�;�����y�]����vP����&��B�S\����~]Q�`ʙ��!WT�ha�䒈%wW��+��)��{|��j�t�h�I8��W��Ko6q�UZ����{مO)B9O(�9��Åc0��,F%��Y�;���;�_pZ���(��+xX�����������
�q@�CV2�f�-YN������p��S	�xj������K�����
�.��;��k�lQ�B���z��������]K`I�$�!��S{f6,����/�o�5g��u�!͊yt�bhb!C^ZU癟~)B���d,����'!w�xg���b*�e}S9�g{��W۲Ф���lַ�� �o�������oY�>�/���:��D���<�y^.��5�B
�Tm
�f�}��P���ޕ���7���l޸��9��._�j�_WGD��{��;N,b'��"�SNϕц'��v��E��㎌W~�pgE�5�2�G9��!VӑIC!^��y��ͳ�Z�f-�
횜1�E�J���]7�����3i��a�h�u�C�>��nof]ؼ��7-�2�u�nr���ݾ&��E���ïӧ9���`+_9�ڝ����@$@ �jk�S���H�D�!�U�҈i��I�!! (eWf�� P>���J/4�_1y���\��F��%���>���B��~��m)>? ���w�12�J�t�]�{��2���=����B ���\��4�('Az�^�M0]�mfX�%&IxL"!�;����|@v�,;+e�1;L�aL=�T+�����w��3���j�G����(���E:�t2�q_y��Pk��wU�����>�˸�3�L��h�����X�q��F��ϡ�S�Զ?6�Y�f	5,R��7�c��M�V�����N���.��N��h�.-��h��w}")(/k��iEO{pO��3סR�=c�Gd.�~�:�=��f�h�!F���_}�>ܭ��k�֜�u���:W[���с1�4���ݕB�r����-}��q�,��ãL������佣>�m��pMUU�ń4km�
lBQQ�r�N(ԁ�c�[��%fH���BP��)?&Z��ㄹ�ښ�$�4�N�{7�U֧tD�t��|O�>!�8A��I�!1�LHC	H�AK �Zk\�g}��� O���T�����B���>�f߭��\^�<DUc�o4��J�EE<������$yw���cq���oϫ?We
�t?�ވ޼>�j�i��<�2�*=~?�nʺ7}G$-��澄�s��_~��$��0$;��=-�@��i�*�����g��_����Mk��o5ߞ������>�'���12�J�uf.�B� �x]H��y x�#�"�)Q���P�AJ���a��[����?xz�V�n���A�E]�b�(�T�,��('�X���DrW�t���yp����J�<���k����gýT~�Qn3�]g`�Ͼ�ɞ��v'����ե��1"�����_.��0Y�/\�ɞ:�3bb����k��/XZ�����W��Ği3�V��u��"%�geb�x�1�9vN��.��&]}�|�[b������NѮ��^�Ќ~�ᚬX\b)�QJ}�N�3��4J`�F'�;��D��UU%b��;�ź]��yl]B�Uk��ުn�2���H&Q � �9�D�")��" �<H$��"�LYT�v��������o>^�$�-H/t���W�.^�<��<�� Q�<�UL�e;H���}ⴎ�VqG��kO�/\��G�]�Kɗ^t ���ۧ�Tp𩝫��<~PW���X~XhA�Lm��yF������[����ߍ@�C�K����ay(F\�BW���w���;W����1��\7UB$)�}y��֍^0��[F��>lg�@�h{2���������Y:'hI�;��l[<�`�8��t��߿g/T��˶�(��:!o�R�.v���oXq�YR�xI����W��!�Z����Y��[����8�AS��Õ���k@�E���-9Jz��[0׸1hZv�����;��PsN�uR9�l=Ѧ�ѐbSh�YOb\���Ef�Z�,�G��R?|`9O%�D�)s�oy> �i�U+VȾy��r���[���Giŗ۴J�/N��^fɆ$�Ci�L$1U&�he$�RR��q������^�7�=��Pk��Mf���}2gN5�Ow=9��y�Ё~c����h5�K:�`��p$��?{�Xf�0c���W��/XZ����n�Q��$T.]� 9g0��ڨ$�PT�����W�.^���=�+Փ�3x���WL���fBf�N^R!�t�2׏������G�!��m�� ߖ'"��AYl�6N���	]�ȟOx��m ���<1�"2V��{�~wwqz��2)��P��;�}~�� ,��7�r�LIA��h�D��N�u�{��J��r�����w_MS�n�C��CE8>����ҳ^�#���
�/������{;13��Ɖ<�S&-$�}����浜�������p��x>�����W�.Du	�֪�]ύ��d!�n�g'����۱j.�b�K��+7��'WH_M�t:��e����q����s���;�4�i��J�� �L*�ku���;޼��0�v�2A<7�,��mF(BAw��,��!`�/k�d��U�YR����(�ZՖ���6�^�jpϺj��7N��Q��^
�1G��߇�q��H@����3Sɍ 9�迪{8ӍT�g��Z1�К��k{��� d�f{ݮ���y�˹�XY׍[t��'dE!l�S{&7���N{��aR��Ĳ���c(S�HK���vSm��``��|�d)���@l9
H[L��6�̶����'�ī���J�8��C��U�k�/&��������O�T���-Ӱ*)�Fl���s���8g>;��/���8�H���tYס`�O�9�hF�kq������I���T�s�����`�)����b#!,���|����sm�(�&A|�m���T�]݋4=,7P���r"�4dm1:����Q��CPĉ��$ƂM�
q����ELg��Y�f�6֠����5#$�]U�{�d���ڮr<�)�[�H���=���r�	�_��k	��e��d�*����e��Yʙ��_�O��Y��Ɂc�� ��߹���!	^@��^�ќM�J3��y�L�y;�_@�~uĭ���{��o�Ôb1�s5ݚ�x�g7=�Y�h�&�����&�ƽ��۷���h��C���𮟊ϳ��	�Ay�^��r8{�m>[o^qq�\��^O�*��)��Օ�&hs�:�3�	���ؼp����z�ngk�s���fq(�L\����j�	��sO�/�q��r��>ɍ�F#9ϬL�Ѭ�O�U�wW��<jՖtG ,Q�2ks���A�/P:Od���QꕭU��6{�3��+�Hl�ٮ����f3��8�����~�2,l~cudI8�Z
�C������
q8��?�yo18C�Okڼ��/:"PZE0^#�N����#x�4�����w�m��6�Udi�A�&Xm��X*��w�މ%�|�X�}R��>�ğG�454����}�n�4%.�n�I�P�؅Bj��W${�C΁��S��v��B̃#)�_]�����.����ł��0Ti!��dxq��|�K�� ���Ҙ�R��,T��Dg�T�9���tk�1R��Ss�Z�;�[���憒7Ҽ�=�*=L��gtjV(�4o�5��7S�*|{�����z���)#��O�3�B�W���{�3�����w�8J9������U�ؤ�ŗ�Qg*gX���&)(�ȩW���{����D���$<7��<�&7�oF��و����kxo�$��}��of�%���cZ5��*j�LW�hqi�6��}Y�5��({�,7�k<LގkƦ(��*sܳ�h�g0T���t�p��x�x!n�<Wa�E���� �&������&�̱���fg�q��I������]N �S�Cp	>���덼���[��������R��6���L�ѝh��X�7O9Ve�+M⣿0���c�ۯ���J�֧�iJ�\������J���Q�>�t;�{}�}��tt��?<k�'F�39��C&�����z�a/ UD�x�i������{��u(�7b��4��r�fP;�u������c�ޗ�ˠ7T0ƙ�5��oF���`�y?x
P��s���	1�4�Z�~4o%�,�h�cɝQY����هEk�`�{�������j;
H]L���fRf�p�$�^7�߾ͼ	eNo[��:��]t��B�pмo��F��}�5�Mtb9����� ̣��_�`ůʪ�./~ va�)�)C��o�=� �֋A�7�Ψ��1���/T[��� �`�l�[�s��x�x�)I�Sa�ao�34DHC }5���7*+/z������q�S�4�T���wbρ��:k�K������B����Re����� ]�B�[�2뚃����Ѹ���ZR
^�͹>�p�y<F��-���&^=U.@3�#�� 0�"l�A�/�V��M�ͫwN2�#o����a��,H��e�I�E7������%�D����ܷJ�BN$���n^�9�2{9��@q�tv���˽/�2��0�q��o�������9Ӽ��`N�)Ěv�i�	L �,�z��/��"�բ1�jF�+X��9`���ǫ��9��|w3t�wkĳ��K���ﶨL3���w�{��sF��6��7b!_0����>�L۸��;��X{�~��>,�\�$�3+$���� ��]�nk�L�v�w�ߗ:�
}t��yv>���k+[-�t]!KDnv_��ə�/�e3)�v��Ӽ}�#*�7sMeP�L�ᡏ�bh��ӽY��V܍cws&\.�jK)��˿WŔ��Ʋ`�c�_!�>��>�9E6����1��Hul�}��C�������KA���d�!�����3�!��/I�}H������4�R� wrPÊ�Sђ�噪��Z�erAH����;J+��!I$����B(�QEQ$QB���cs�$�����I��[��舛��������������==,ɑ�������[@9m��-��Ns����s&L� >�9m�����^[@��@""rppYɮnYe�����}�G���$/"��)��L��7�BKH�@a�M�i�1"22�"�2B�QDLQE�*6A��TffJF&��CN��F$E�Ð8�E�JI�R�y�_�<��K�ET�B���g�e�0����6�6�M4Y�^rד�z�CL�!��i�R�cyhѳy�mEM��I�sy�H*F�(�Q4jҊ�E�C#* ������'a�	11�#	&�PF!�I�ryK��n�BC�8C>͒ų��j�>f�>�h�r,�F��7Y�n�A�S2w	�����ѥe䛢��z��o{;+�+ݡZ���(Wd�,��zQ�]�L0rԌUV;l��|��ɩPG:
݇tq�Oi��q�*�_�^��z��ؙx�P��w���ݘ���Y�揮��bӾ�����F>�6(.�D�u��j�o9�"��ĩ�Z!Ay�ոP%壆��9Y��c,q�j�dd`�G��Y7F��Ɋ�%zp��#ID�`�7����O����z�Z�H�\�|1OP;���_=�Ƿ6-{:2+.t�hP�3���͗�͔�b.�3����1�% ���~Y�4#ph�>K>�#���˔�y"�;Ɗ�W�g����Ē�$ �:l�e8��m¯�=us)�'7ܱ�� ��+$M�p�P*4˔{�|�<L��FH�uAbL�j�*���
��T|Q��,,��~���|o���#6^�sk<7���`j�鐖n�T�",��Dhue$�">ޮI[�ux",��Zp�f��!*���l��e�R�t�A� hAx���&���"���Y�tҠ՛�]�;�N�x݃�h=�Sٴ��6��Ʊj(�������W�)�l�4`�U#�\f,����3v����(+AN[�^'5]ɜ�����x �(�>KZ�,kMٽ�Ρ���Lٯj�v�	��tj��n��L��]��1FK�S,��J��O4ᙜ�u�[OMq�h��gK�l
v��G��Yʵ�&��Eb�H�i%�qƮR�MW/v�-cj��q͞��W�t���ܫx�����+�#l�����g
�ɞ��}�7��mu��;�34��I��%-��6Aܮ�=۱}S�V���Vߎ��^�2�1�M��;����O9��{��L��MQ�c~��ٹ��r�r�kt~C�6iM��9�>Z���xKf�h^dL�+�8�v���82��٭֋������.Յ��Ĉ�� t���|RÀ�,?�_Z�L��_n�M�V��9dmҩ�$Tw�[b� g,q[��d�gCc0,��/5��s!M0X����2/[R�7��� #��&�V���iyy�7Y�w��b�1�+��*"��к�4/l��Q��=��y�"F�����E=�z�)�%�g^�]�p�qS��p���� ��-�\7�|�����5L�B$/c�<0i�4�|6s
x�3D@t�2�Y�A���Y���S�{M!7~{��r�<�e�5E�>b7yq�7 �ƚ��Ǚ��LQ�
��t�2n�P��@��]�����V����rBT1��q���$"��μ�'P,8�����9(ؐ�`���,p�P�Q�":�'p���˾��(�t'���h�嘲��a-�*�P�������&���ۖ��2҈j��g�W>��|m`�)������D8|�w��z�F;��`�y:hЃ$�xR�Rϵ������e�r[�j�ւ��'�EϪ�,^O��oB� G��҇ÈD|7Pt�x\�'�8�� ȅ'o-���y��a�Gc�kn�h^dNLj�#;�L�ѝ}!���^9��fe�j�L��5h[;xְw@r�vDR� 7#�W]���5�Љ�
ד�,;@���쉷`;�qW��T�W|�2�P��ϝA��4�b�7!�(�ֵq��^��kX�γ3�ktS�{ۼhΪ?�0q�I���#N�{"�z/B�pм-�zE0[�*�z��9�Y�Cݠ3���)	9���O��x3y�0)������]ֹn�Y�Ii:��@G;g�4ҲH?%�����4hKD"��$�TˁI�9�[��r���_U
�4�M��m+9���GL�իp�4\A��RWb����7uN5�g	0ì%$�-�m-&ܲ
��P�Xgk[ʕ�r��v��T}�	}�>��M~UWq���2����5N��q�Վ�sd4��r�a%$&ݣB:Àκ��3v��
��Ut�ބ�Eb��ߺ�������K3�|!d���'�ЈcĆ�s���oP]x�`�����;P�r�,{�B�N�sK����M��N3N5w�c�Tca��~&��V��E�>�L{��{r�D�� D3�	�v_;,��-2��� K�	s/�z����λ�m�w��4"KRn9���k��WN�Z�^|}�xt��ț�;iÓl�4�h�r��DL�cn:����K���Xk����Ck� C)	:V{3
�ᶱ��'��ȵ�F<��q&�6��*�T6⾥���7���4%OzI	f=+m��i�a�UsIn��cc!�"��Q;�7�<d����q��AH�*��d�E��@Y�˽�7i�YW����N�Y���:����Jݨ��B�f���hx4|﷬�]&��zޅ]G9"�*]*#��S�D�\��H-/4�:'��c	��#����aj���6�x\������u��P��]���k��;�\�	��ۃl!�%Ji�w
�}�U�uU�$���)��p�ǂH%i�Ӧ.�5�]'���7��J��٪��[tAۋK�zNS6#K�f_WV�;8���ݦ�b%�*n�J!̅���U�Q+�]O��ָ�D�mO����Y-i�Ԫ0p�NvL�(~1�]�Y^'k�M�U^M�ۍ�e�Q��A[D@"�����3&��[�K���]D����H���n�勋�H;zP:��^�s�:j>�ׅ1�nhY$ �4q�)�zc%pv�x�����o�A�l5co痨f��/���;'�pǆ�K`Iǣ���x��E��������%�Sa�mք���>����H�l�Hd1���1��aɊ=j e�J�LᏵ�'�B����>�T�_T7�!D�>g��v�.�]3�a���)��cc�ii�����!���Pۙj��ի������q�5b.�r� �M����]j8/;���F{�rp���m�,4�Ą����.7��Foh�3�;��keV+Y���C�O߽�^��1��I�����߳���1�g.uX�Q�b�~	�Q�귯l9�."�Y�2�ٗT~Q��T�+5�(+��7��:�$�zO>ڪ�����P�TTI�i��6����M�Mّ�"���!(H�""-D�	�Q?|�{	���h��;$����bc��\�
i��5�0Y	%3'f�m����1Lލ2�e�SAc�ڨ���	����.���)X+�{�� �q6�.��(V�5���?{���g�GG�C�\��V�Ϯ�2Z��/Y���׳��vg�źg���'q"W:i\ք\]�c[���V�J����Y��#=OG"����F�?쪝{��\=�K6؍�n.�]L3cIs�m�Lp���;	Q}\���J�b�I�/��pU��~};L�]&�g@�?�spj��9�\{�Sof��Eϥ�e5�-�ʪ�s���;f���i�ԘA����D�a�Am</k��QqQ�k�AP���{B+�[b2ld2�Wq�L�g���a�G�R�(-�N�Ί�$ͫb_K�����y5u�"-�T�*BR���y�&9F�	����7��+U��<��LF�dUPă�ݹ|h�����UT��4�	�>��@�����9d�Rh��8��Z�;���	�!�s�����{m��� �\$�����Ou%�4�����|sbۖ3���%ʆ�L�������B��5�q��7/R�O�k���F�<��޸[��jŸ��E
�"������^.n_�&�[�������=-��<VD���x{�=S��^�C�x�ne�Uv�E���k]�r����,U����E�ݤF7�d�Cy���(�'M���9����r֐���J���t7fe�#!��K�+ݟ8�7�����k[h���T����6'[��v�c���
BN����1�?S*���|�Dim�w;��^D�V�nV��Z��ߵ�s�����` lV���$x	$yoTЇ��u��y����vp9[�8�ƨ���vV�X�qk;0P�(�1�vj74�̎���ĳ�D��ST��M��@��MW��ׯ���X�yt�ϻ3�(��b��DIL����7��v�>)T�e�S��^.�h2�x�1m\<!��s����g�	�!�s��� �e- 6Ѭ~O�j����OCDO�dh��7�݃l^`((&K3�Xa��~���$�P�)�Ar�2eW�t�3g��B�F��e�����'O�wn��F�<l𧇄�b��wr"Fܑ���)�i��'�-�� ����������~ƽQK"^e��@���*]�����a������c8�����b�c�U��5�ƕx�L+{O��4c
},5-�����RLO9��<V�z������C᷽�Aa���N5]�rS��@�C���Z�����\E_W*�S<{�16��f�i���p�Ҽ=�!B�yl����}��Ü���X��&��~�B�Y�*��v������x�E����FO���
�&^��5"p+�����΢O{�j�V�\EB C�n����=3�b�G�FN�ڟ��]Ϙ�[��'��厢:艱�X�$�xE��~���7s��n�^k�Z�\��T��x�ӽ�L�k�d�#�!���>�ޒ
���;�HE�n�;�(�j�O�tp��7��w�� 5�k�7�Z��<hb^ 6�}��� \ؙdՙ }��y�7���g�2�ɩ����MD\q��$��C{��S�.���{5�b�wYX�o}����c�_2{� E$��zJ(��|�J��'� m��%� G7UW5V��.�,o���j �8�@Sq�Y���iղ��H�,Ċ����f@Y��,���ͱB�OL�|�Uol�LT=�������\�vӑ
gY��0�mc����@��YNK~�~�{ywM���m{����ƶ(;*��E�Y�w����lK̠3s�%��W���0�jrS�����]G���ڡ:f��������g7;y�Ę/�ʻ!wU�]�W/3�v�q�-b��G��Km>`xxi��ǻ�<����;K�c2�3{��z "%���g�t��}�J�{����
���!K���q�~u��3G��wU���p�xE��y��]����~����J�Fɛg���*�n��pB�U�0�$�Dܟ�|�4|��2�ĥ:��9���b�P�j�Y��/3��$��o @ѿ{h.��l>@��|��:�DC̵ƾ��< Kl@�s�T�JOe\��a+u��-�m�u!���qX��efA�n���U�w�i���n�e�9k{v)��F��9
����̛����"��RM!2`�v�|x��~��k�пQ�9#O���z�>�o]�6�h�➽�dz���,�T��w;�%��śc��N�n��k�D���[*:WBo^Ky��W��ӷ�zr�OY���� �r�]� �}�|�hf����[��Uw��h��T��P��,W������aJ�ݗ�W_=�>7�D���]���DB<���4c���ۛr��Ψ�W�ϖQ��c]���/�%��%�*�6�G-y"�@�}����v��Plb���s|f�&7pf�H�u��KUN#r����d�i�۵b��#�W&�e�E��B=�G8�t�hs��:�o�iCJ�q��P���d��7�P.ˎ�%�n�JH,J2�`�$,X�tOL�:��~ ����߹9,��D�����2�\�M�������w��陙����5bnn&�"{��,�����z���г��0�{ {ޯ��$�I ���"I�{4���o{P�@�b|B2�l�Y�SL���9	�O6ܐ�%�D�)�0�I�6�l8diHcj9v��%d��U+��Z2��ӥ�!2�ӵn\�$eή��b+�đ�-�����8t眳�֝'��"�2i�$	���_8R�ьc)3#�n�$�A��n����PE����F���O^��UK�\�Gݫr���U�^�3��^�u:���֥��q��m�Rǁ�ȁ����3�D)pw��R��Y��l��9�&�����٧��̚��NuE���z&�#�:&�R�z�ˢ���"��nmvrzc��;�����{}�Y�yjjʠ�	u|��	��	��^�;gv����������K���_u��
��)�+��8��\�6�h�˙TꙢ��uEXp�'l^άX��^<�X���y�,�2^���u���es��{8�*S���h�n{(�ui�RU�B������qv�f�;5�Q�����q:����o6��Gv�f��U�j��9[���;*�w���_#���G�z��I�o�X\�n����$M� V�gLH��,�y՚D`w ꬂ�$�2 L:F�>�H��Eꩪ��z�)d���$'y`s�5�+��`�V���`�߱��j�"��Zʣ[�9��Da��N�sSFQ殯�㜎��#R���n��\�Yv��(�����Z�n�/cyhZ9R��V��jU	
�M*���7��r�ʺYN�J����G�  ��a��A��-�ї��Z+iv�˞�Ĳu�\X���=���ܒ��m�����N��$��L͙�3UD,v�ڝ�3 M:V�������f�ʧmF�����QDݢ���$�Q�X/Yv�,�aWQ�j�P�$���֌zľ���ԺG�2>���A4�.&9Cq�$m"!�$�Z]6��O�g�LA{���J��G��.��Z�HZ�Q�s48�K�����Z͗�ѥɌ�m"C�z����Y"�4h%z�еZ|�f$nHa�����>�hP(�N�d�/D� �wT�ӡx�����Vr��倄%o�u�x������Ԕ�II����G�>�ҢU,�q�윿�:�l�}4n!���/bWW<��u15�{a�x�ݯ:�ni��\����-�٥�{��'�i��qh��Dp.��=�@`�M��4ʭ$�E�>�LzZ�w����"�x��j��������L��HSj�w� �F2)nw7X�%lI�v!��4�8>ɔ{�<��C:�3V)��+��_��vfXj�d�a��@]g�ly�Ҹ�9rg�K����}�? 9���R�9�H�c������VbO��S� 2cMgl�Cw�z���˛�JA4�(�իr�{-V�@����OR�%�uM�Qe��^����&�[_^U��9�]A��GU[�����	��:��w���M/�Xy}���-fˮ�5�+M
\:)��ᚧk�U�sR��rO*�tݐ6=�"��T����t� �vJ.�J� �M���[j8xg�t^gJ�g�1�S��m�$h�'��*o�o�������t��C�;Cٸd��$�g���W��I�?z?	z��G'"����&�)EϷ+���G�o��0���ÈK3Z�{�(�u��qH��D9w��cϼ N(���Zy�{YS��5UQ)�׭��#�dKw��mԤgG�\C�D	S)�ݜM��v3�=ݙ}$����z;�vݚi���
R7(3���
��&�S��k���\�n���W����14�Q��~���F��.�ξݻ5A}7k�M�F��wϢ�l�"��B}�;�H(�7��8�"�[�Sv2�c��*�q7��-6�!˵�v5�]l�ju�{�\��BKS�&�.u��ਸ����L�̗V�h�<�[{`����gQ%�l�tS��6�Ʃ���4%Oa!���XV˵(�ժ"Jg=�w�F�͂��g�t��N�-X��A����^��@��? 
�F
	����za��N��N�<HL�K�V������wzt��4�i<4=�E@�0�F���=����p���n�5=(����41;���r��޶�hĹc�ڨ�ѼO�p��]oGT�W'��$C�x�Q���m,�x!�%V��=�al[LyNkDx�x�����| GHZ���aɚ:d'E@h!^��#��+�9U������$�F�ʕ��5�̡�PK�0@�C+%��UU
�wwbƌhiȣ-��j'��J"�i%N8�e���(�S)�>N����Ӊ���Xک!�ٴ-�s����s$:�z�H� �E�r��,�eFo��(��)�V��\Ԩ^����������A��tCph�{�"�D/cFMD��g�x0;w�� ۬�	`J�[�yd����V���li.|�v|�&�d^��z�TG�
C](aO����>N���u����I���1O�#�ѓ��g�6����X�>��ML>�j�%3��zc�]t�p;�V9�q</6j�P.*4��L�?
d=�#��gS<PL�K�n_IFR�=������=��Y��f�B��;l����,���ۼ��[��<�����1=�<hb^ c��"�,ܷUz1�Tʹf;,�����672��A�C!k6��9��J�f�v�fha�����X4���pk��gu]��@B�I.���4��A�¢��P#i�f)YĚl���Z�X�+p٪���@��ִp^%�[V���H��HT%��/��)�7_��{�4:6}�9��7���g�<=���U�x��s!��+��u^�ڼ/����y��{�nZp�����^K�f�/�M��l�՞ĪUd)�ڸ.�u��+�#^�P��<�^�����lH��tE���%�S*<":��~���m�f��������Zb�D��z��SǸ^���ػld�4f�>�����#����HHRC��b���}4�z�:y�˛�D�{���fS9#z�'�۽ፗ�)�TD��`:a�`����	����<ʚ^��z�-�r��L[T�i�s�a�C&3�M	k�97���l���3;"�_}�ƟEj�w��4`���m�����^��.K�s�"KB|.��k��E�v���M�.��m;�غmJ��~�=t�(��5�n��}	�!�s�� �e$�Ѽ<��c��~�4�n�v��B��;l�!��/���zG{�1�[������_h�L�B*N�.�9�������R��)]�������?����q�O{��%D�lO��$.�OnX����D�Q]�G��f��X�/%϶��/%L0��~��,8�g���>[��-���fݜb��1��B�ot�:�� 7�}��#\U���i�.����2f�囖{�&��=לER�:n$�.��	��{�����
���:�#EYc�}�g�f$���w�8@�n�UK/K6����Wo�C��O�hv��\v�z�_!�O�tH)'����._��8�����n��jw	��h[�8��6��;0{��y)m�B��͆R���M��5Vw���I����s=y޻����-a�JcGP�b(-� g�m��`:a����6�sۻS�@���^赜�m��ի�+���r�&��"�c��6��F���3>s���xq'�o,�+q#*���VW^� j��[N[��K˯�񯳷�sE�q��\���r|�~������{E��g)!�������s�� ��w$��� _��<-M�`�E��C�f%_�xx[i���<c�`���g��7�<#�~����Sݏ%Ϸp����^�=�m�˷{���gFw7{���<6�[F=j�^֍����'s�ķ%p��K��f�Sp���(+ߥ����X��d;'ΘZe�&]�݋�X�@���g�!K�;��A�(Z���)��qEpD�IB�nsSs�Ѹ�I!��"`��e9�)���]vSo�7�qQ�^�uo�7P��6�C����$#��C-�J�Kr��;���o�9ʽ��(A�:9�Y�r鿝�{�����	�Y�:Y�W���n���VbMĞ�
B�(�x��*��ڊ���n��e�CD�>g��u]&�g@�>������������z;��s�.���C覭]��h\��SQ��,�4�x^��Vc���^>A���()�6�v��Bf�bx �{&�f�  ��� ��N�"ޡ=>T�,����kX�w�l{Ël����]���Jg�&~��a�n]O~���-�m��M�J2|���DM p��Ėl@�I�@������Y�۪Y)�[�o(;@½�o��+��'c���-�
X.�l��T�c*W}�����(�4>��{i'�ґ7��B��M��p�QD�u{2�v�Ep_Dj���i�!jn]]4��A�����S��*8f��+V��q�WwЉG���!��EKB���ы��IL�
��@�,��x"Ҥfv���o��U��f��E9���rO?�߲���Ͽ8�1��Q$-�ڸ.�w��궪V?6�<w�M�}��w?kxѿVp� ww�b�w� �T��������ly.}��>B;�e�ƻth�� t�I�P�&at�9�Ƌ�����Wvxz���e��K��,������o��^�� ʛ{&Mz�U�ĳ���$�^�ghG�F Q��g�6�Wz�X�m����li�A}������4b(��$�g����c��O[DHd�K�e^����V�����\mp��E>B��sn��'e��GAP�Anf�-<.�-��[�\D�[����m��Z���=)��D�4mΨ�V0X�Z�Q��ټ�gWgr7��솖Jk�م���[iǙZ�m$E��&��[�y�p�L��(a�hax�L�(K``L����a/��㝾W�a��q���5i��r�3��+�� �.R�cH��f�*"j��m�����p������w
�я(;;��1�jS��"e[���_�V3�
wZ#�dDĞ����:����v��C
k�����v3��\w�)$B��Z\��i��9��B�z٦�X��΢���]�2I&�@s��6{���	c6�w�jy.}��>aK �=q䵬 �#z4�(p�0��P�}e���u����t���)US:5��y\t�w�.�u�yw���,�#^a�Lh��QS9�����jT����a���U-�<���V��d���m���i�!L���jZmꠗ�X,�0�jC;� ��S<ri�%j��b;i��:T����,���`UV�aز
VC�J�J�Htm���{J"4���p�3�>m�����@NW�\@q-j�Z�XM]>JPk��"[Y�usI��P��j{�5��K�۽7��d����5�,�\���x������k���v[�qo�}��K��dU�_]ƾ\��4���m(�
�jnⒹu�k�㌛;\�]ηgr���j��Ǳm��0
AZw;�Ž��k��iR��Ηb$M_:\p�U�X�{�#6������%�D�>�~`�b{���:�飸K�&�\R
�9A}Y	���T�t�%��u�4��\zm�}�X�fKX���Hg�6�rM3h�i�S���PPX�K��6�2�l�h��,5�tQL�n�+��W��5��]M���֮�~�C�6&r���&w�Q��np;k�>B�d������#!��T}�w&�^a���A--�H_-4fq����Y>8�K�Q6�f�DHۑ���(�1i0�9}�{���?w�������hD������������2"&D Y�Y�&L����;;;;9�h �-���������������2� ��嶏M�y�/-�m��ss��8,��Ye��>D�-޽.�;=�68�!i��MI)�n$K	��P"&,��$9�-�LQ2�e��QELH2LED�/!M���[��QD�1��jI��apH\�Ԝ.�6�ߣ�:-��h�1^�AO!T��(���u�s7��2��0���c�ˣr���J�>)�#)E�<c��ALTK\bSM�
P4�n"�R�j��ṁmy �$9��2�'�)q����ZH�	�q�qv��,9;p`��e�]ȷZ��3�{��yhu9���ɭ�}U��ݡW�_q}�Y�Tgp]B�b�=��&��FěAmuAToxaZ�{��(R��r����4q���]���[�ٶ_*�]8&t�+���]:ol�|V�RyG�d�ռ�Ү�[0Jё�/��zforؚ	XMɞ�4���N�0������N���+��ܸd�z�[������Ӗ-������ֆ�}����eL����7�9X��b�jq%]��muX�H����Â���oRk���<�w�նی0�-�յ�Y��Ww�iZ��[�qggu�{ս�p����)5�6����HC��C2Jt�=v�^<�{,dV����b~�Ts<��.�YM�Q�7���gH4�q��{-��^�n֭�������DK<�v�';-W#��%V�?F�IB�&J�`���,KWY�C��ev�WA��S͐���l��E8����y����iڭm��s}��2g���$��j�*�f8�HP�3�Q�[c��a�(u�9��[Θ�N9�p�W���X�^�,f��k�q�rQL�Wi�(��r^1�����j��f�	� #3��`(CQQy�&ش����)��>i<
�e�twBCZ�V�<��~,��z=�a�'r�T�Q��廥jzw��W2q��g�Z�b�,jPѷ\{;=��b��q$V�7a�r�-�8��!�
�{�����p��{��})]�o5I�MwL���v��f��t���]\]vgSW�.�w�1P��t|
N�dL�bɔR,)�jC���P��Z[3Ul�
�1;9O���d��R���i���[�3l��~�\�^4�D`d�K�u^I�)h�m�����
J��aDl�O�dh��6}�Of�w�ă��&1t۽�Յݥ�bw�&x���@Z���[����	�Yߥ��{�p��3Z)
���M�B���1V�6�p���yB�;T{b-�O0[x	j���������,�h���\�o]��w��b��덏l�Ӭ��	׻.�q;�k�#�pR�l���/��챜�1�p�������$�ĺ�G�T�3��>���0���!��s'Vm��R�lo������Eb)vv@��{۹5��N�˃j�g/�>u�U��Z�M�[kc��iP�]݈�Խ�:�$� �8'*��52��Dc�cq4�m7~.$�� ��4RȐ)#'�HbH�&bHf��p��+�;��ɹ�<�[6�V��ku���0� ʫ��LPi����(������ �8�	�7AL��-�egYw���YW��!҆����3�k:�<����I2PrH��i�� ����q��>�ף�o5>2�=�U����k������c��DIL���8�<-�v�gq~�-���ii�7J0�iSl�W{�;��*���uĺ^���(�N�#zM��iܓ������S5�>5�v���iM<��۝��6�oɞ41u-�b���D��e�Vd,��F�[F!�c�2��浪�]�&���{&=z��J�X�Si���mO��$.F��'A�-(��kK�� F3ux�������F.UQU�v��þ����~����дYX�Y�}R��y�I��}�^����۰���|0�tcm���hF?U^u����a.\��9�rc��M�R���֗�;ƳF�
��c"W�t�9�T�(2�Nm�5Tu��D>�D �i ���T��3A˄b%J�D2L$��!) LH$��g���'UԾ�˩�z4�s(�o� ��YL�g5+��Жz����C�ݘ���7x����l�DL3ch�%��� L�_=ߐ��� d�I�]�Q�3-�7����[�b�A��8}&}�ğ��`��7�;���0_��^����ݮ?A�r!�w�o+y����вt�s�Yi�m��i�_�;�>�{2`KR5��%�p4�!�p�`!�QLJ�J3#��χ���4��Vz�}�5U�d(b���RF[A5�s�L{���l؟Bȱ;h��ҚJ�=���n�9�<�~O~��UCZ��I�ͣ�{�UM�G���p�q@{����!�Ě��Pkqfm�1�W�)�{͏���W���>	D�Y���k�_��)�Nի��{\[����7\�"���}��P;7sPne� �D�.M��A$|��H��L��^M+7d�ꏞ\}�s� ��d8���7Y�ِ�yC�=�|�ѿIW��ǵཀྵXѾ��^2*N��-��\�����~S��}��1r�Z�c_ژ��p����0�V-�]����`�ؒ1�TB�}٦����G��X�B�$C<Pu�n��5�y�li.}�𮻡w�*"��1�n���m�^B&��=L�)`5v�Ǣ�<1�P?�g��Z'��B�OşI{�ğ[�ɽ�k;g��!z�/���-�2�ڔ>�k�����H��d�`:L)���6�ݑ��p�n��˗0Ͳg��CN��2D֝�2#��y�\D��Y�XB����4�&��ƪ"(���w]�z��7w~�ç3�I��������S���Z�N���uK�5D��B�Z��mv���ף���X�H�
��DSdRqxˑr���[�ۼ�xv׳���l��Kr*J/��-����<0H&��~1���-�,�"S�"�Ut�(�@�GP�SqeY-.X�/z�Ro��� �]�"��aP�_3]竀E蟟ԶԃB���9+9W������vĆ��\��I��UT_�~�,����Y1/��˝f5�^��aM%B��{J�ݗc:�xGofvt��#��׭Q��f�Ej�=�M#vF�g^��5mb�a��K�knϘGxy�|O��Pf�kԮ��
�r5�Vxx;�7v�7�i��ճ���6K:)��!���e�[� ���6#�
d*��J,��Yx��" ,]�x�"�n Ӝ-��M\j8�8gw,�^ �oN33�UW
����X���֦P�6R'm�n�Ԇ�We:I[ϡ,#=!i8[fFK~�7�[4��d#KZ�V�;ҡڭ�%_�Dc���W#��N�#[�1nc��I���ܯz��V�Hҽ)�8�m����>��7���?!
m"�	ƔnH�M |-+����/[�+0&m@��H�Sk矫��e���Ĳ���N��2D���~�k̙݌: ���I�Ds�'�ڔ���N���{#����'�����U�54%|!�^��e�S��t"��5f[AMe�-����}� N����d"�P���{8]����x ,=D����ǽ�*ų�V���c]�u�_�;ݾ���>�b��rbu�;�M��v3��k\p�ݽִ�
(�xz�;^��呔�'U�#��M���u4��k��	����~�G�j�$��k�h3�S9ۨk�Q�Y��{���y�V+>�i Ʈ�ʉ[SV�40��0���.�.<��y����\i8�l��;�̾\��6�4�P�rܬt�Y����W�v�I��V;����\�*4��u~�A�a�l �DB��[zL=��3^(��c�	�e�ba��K�n>ϐ����������P�z崝�L�L�ӍfO��5�G{��}��hx�eS:)��!͓:��3ۛ�}�@J�h���E5j��Y�\�:��7��8��Ͷ��cM�ڍc<�{j���fDYR<pY<�&C'�������FR�xd�nf�R��^��{���Sۘ�B��;h \���;��%n�!���w�~���c[S@�N���aDe/�O � Ai�7�-�GO�>�����Q6�
w��r5t��fB��gz�&=��Jy�؟�hP�`�w��5�i����zB!ggַ�>�Y"�m�`�ݯ��6aa������<���6�BQ��[�g`=���H�f�/$C!u{@�
�]=8��Ri�y��3w8ֶɠ�+��6)D7�]ˢt�ʫ���z�F���<U�K�u��v�ëF��7�pE��)ަ%��1��H?;�#^�p�G�Z����֑]�H��6D�3[+<"&�;�O���f����k���Z�@�z����α�{�z�;*�dD=��I���Vz�gQ��F�L�	�C�xO������Ecd�=��Ÿ ^�2,��U[���ծء�S^�UP-���Z����&�v���t�תbΘNt�4������Z��!�u6�{�HeX:^꼂2�c��w��#��4�>�IP}oE�Y�
���u�0@]>Q>��� n�E�f��2�R����������Q��4%�c�B�m��ۂ5�+C��W�q^���\۸_W3�ӂ�=u�{}O�d
M�ٍ��Yk#t�wM�y6��(�(�1�LP�P��t��V�fP�=�i�L�M�0�2��*�is��Rw�t����O�f9F�Z���6�
e;�f�xX�)�4�=�͈S;��\D�a)t^��!~���m�ϭ��C�NA)@h������ٞ+"%ĺ�^�	h�*�w�Co3��#���m/�Ǽ=�iR_h���1�$�z���6�xt���@��G���T��&�����^u¹�U{I3�k����� .�w�nY�y���+iw�8*�v�7�����8Im ��=hk���D�Z���dX���&����T?:�T�E�y��i,j4.0ت+h�l�ւ�(�LW��mgֵ���!^]]c�?]�����q�Nվ��7Z
�5W���mK�l=��bUVUU
ƅW�`c^���$�N���i7#��2INC"�! T��9�]Kf6Z)�aO"r&SR$c�5��&#I��Fo��㹧���S�g���WQ"��#R
4�okJr��5P�:�������鵥�-4�[x�[�[٬��{E��d�e��7�^��� tM�Lsu(�P��9	���w�,fI���R�X��
����_��@U�ۡW��|+�n�2:ր�%2
�"���E#'ϙ����Tn��øm���L�sZ�cn�=ƨ�5�f��� N5:R�L̤Sn<u�Q
��=R'B�w�{ç�Ov@�^��a-%:�H�鷸.����.��n�F�WFEj�^[T�8a�|f�=]l�H�x4f�kZե�����V�A6,��
H�?(�� ���GZkf��z�ԝ�Jދ8ߥ���8�u�	z�BS�L3�X�$8��i���Kt��sUn�,�f�#ݪZ1�!���"|@"$٬&h�p�5����G�o6fNc���m6��"�>@g�_P��ö�VZ��/&��'DQ�a���8��V���ԫ��0� �{)r��vY��Ρ��z� '^b<(�ñ/��kg�Skq-!��a��@�u�HC-2��q��K��\m�-m��qU|���=sp�Ĺm�v�oR���I���j����s8��Z�Л���k��.Hi���\�Y;~�3q�V]��i��C�n�X�P��S�&C$7_*D.���E9�PhP��Y8��S:�'F��w�z�\%s-�`�ݪL�Ε�*���R�1��tS�q=��u�$�	-7}���Q;�ܣc�r3�D��6wDN�ut������}}��jWw]��d�������\n6�rf���{�.]ݼ��>��Q��q�T�%�}���j�'�T�C	862�׼b�e`�8�h��k��k&`Y�-�!</�HP	Z��:���S��!��:偖[E�@<�!����O>HUPHS�P�i!iOR���ݠMC�gU'\�IIi8�)�aL��L2a��M&Y�0�l,:��V�J>D���4�ϼ��)#�/hq�g r�C,�����'P�V-h$T��$18p�G.�v�I#����C@~G�ӓ��,DKo��6 ���-�����5>jn{������ze�Y,Ȉ���{�fff�{wA;���f���o{� w���� 	��Z���q����T&�]�v\H(B�,����B^>! ��3��rBd����iS4(8�%�$�	#p��*@��6V\��1�$AO�N�nL+≠K�TLEҥ$SX#Ϯ�_��=B�$���{�;k:a!6ժ��ᯥ�:N% �)&��bO%@�u:10Uj�Ud��#7�ݴ��#n�I��ʒ1.2��ѝ�����G\��A�T,�fh�mh���s���m��[�ë^u�RB����#.�����b%�zioX�앷�1��̕�:�͋������FWH{w8�9��v�SZ�V]����"��k;�����u4r�:ƫ����}1���GA�ڛ#.Đ��N�x��YA_����A��kƟh}��Gq��k!V:��L�nK�N�$�׍h�<wQ�5X`T��_K�_}�������k0(���oNͭ�O�c�8���M��5q�����@�d�j��\P6��Qε�N%��s4�=�*�c*¡uou98�T+37S�oU�&�j�{:��Ґ������⣈ot��%���3���D�FIp��C��ې2�t�*�%d��Z��]*�ר䒛��#j�M�P�Rf���H���y)�5�4�<�cȈn�u#�2���>uM�8fLr��Ӷ-".�B#×GB�>M#o�p�}�x�ni����E
�v.��$�s,e�٬G7j=��iηld׮�I�'�eP0�Gl�O�,ح��U���S��[O]�W��<
	�:�$��".�D"v���4��w/��a�j�$4�k�(/��K�`�{]�	�w�r�����J�I��f��J�V����O�1�R�"�Q+�#�$���s�d9��Vщ�v˔J
���{������pٛB���qeE6qƠ �Ɂ��M6\b'}G��9���;�%��BZ!�8�E��&TI����v�v��*��E�A�Ҡx)�g-�#hvFV�M�W�<��}s���m���ܻ%��}#M�a1D؇Ȃ�p�C㵋Tp�.�mgu?�=�3�U���1kS�/g��x���|���Y�QD��MO���5�Vk�xSҕ�ׇ�@*qI����Χ����f8z^w/ � y�����%�l4ִ��)�8�{�7�M�l���M/e�A
*�6��E�P�-��O�x8����P��H���A�iM.�#S ��f��S�5ilr�D��4�M�ҊB���u��Y�!�vS
,�� ,�	�xY)�,b"�P�w��c�����S	��H���g]e��	�Y�CV<e�Q
�9�]�u��CX3�b�@�}����95Y͚�l�<ں.�u:�;1�jS��ڦ�C7t���������z
���Lo���}_f|�>���UͧcBT��H�K3����}�T�T���oL��e���z�Ƒ��7��5��r���ƨ�+Ĉ��z�@ �IQ���bgwd�{n�ْE=b�^O�T�+q�{�nCӵ��.��%�a��f�V!�Iƒ��ul�G{�%�O��mf��z����J]q�tCh�<<a�9ew`�蚙L�%阽Ӑ�oΡl� �����f�� :��,G���*�o�L�կ��=wb�WiEQ�S�?��5%�=�k�UK��|t�܇�����h�N�i��x�xS�����L�O�����y���ݏ�	���;��JO�\蝎�z\���@nƖh<���aw�����2��Kir�ћԢ��|I��h��qS��>��tv-�"�OF}��m�9-��֚Iw؏���M!�XY;�!�3~KY��Zk���x�9�i�[�q��qv�v�]���"��Ma���� �#�u
L��Y�e�)3X�BN�>%�zԡs��=߇�5����Іw��ȇ�`�����L�?nj�c�=U��
�Z#�cĸ���z+YE O�y�SDP���	��.�u;�k� p���
2	�1w�Э��R��c�Y�H�� ?!(��w��:w���N=�D膸'K�-;�拤����=q�y[��*��
V�(j!�[��5�G{�����e6�Zes+�rOc�!��<��%�n� �.��>��x�i�SV��P-��:��v�>;�jr%�TB��r�f�BT��~ C������i�L�O��G]��)3��I�]��ł3��y�,�,jq�#�э�E��X���<q��n|�د���p�@���O�����w�t�J�e�K��j1�-8ݱ�/�(eS��c%��QSeic�6�}���\V4�֦�<�F�ʝ����ң��f�'Kd��[��()	�Dvᾘ�m1S���S��i2�Զ��V���pn���1 ˸NY;��~�+�h'��U�O�I�yK7��~��p�w��Wu�`���t��3Z)
�8�	��S����Q�0㙐�yB��6��I�Sf<w��.����?6*rm�G���q,����Z;��.]���q���@�N��v3��k\I�k���M68�l���o"� �l�l�S�V!�����7�p���m�9�U��(�M���oU��c����aV��t^����Df�(����̪�L���)����n�)���1�g^��1\�xˈT��^:�G��+[�5�;b����$�T��U��tkM��Kw㚯K�)A�a�'�$���k��84P�U�ݤ��r$�	�F��K{���zq:�&Y��XH���C/�0`�õx�j�+����<����[S4����uTA��HE���iIid�`�Y�1�t�l��eԦ\]?M��陀�hĘ��#�����;��r�{t��|bp��{i�5���[��&���`�[�(�P��;�{����JY�S˘�B��=h��Қ8y�к]�ݝ�T�e�dh9�1���d�O "(L�l�VCoZ�B��'�m��g���
0�Z�CkJ��TL{�5��R!�:�(��7 `I"d5���`�54����^K^%Ĳ�f�	x�*!���p A$��1�g��ژ}�3E�Fy;�׹��Z�'ͮ X�5�;�t/��H�-!n�]�օz�ϱ�gW]ŲI�Ki- |�>ߵ�W�!�xx_�\s$�zƌ���×#��\/�����PN�:��Ą�۝��b���WjR��CtbK&gof_S�L��,X3j�t�C�i�%�^:1��{�|Ꙫ���8��$��m� P�#�$--�*H��/3���y���oUߔm&�h|��[K�A��ӛ��R�Pf��*�Q��$���w�Xh�G,z��xB��q�:�l�S�p\���Tz%�l�E�a�NF4ڍ��#l�v�tp}��,��çn�:{ip�>�Y���
r�����f4b��ϼ�Q꠆���3�p�.6O	|.(��oTs[6{�e	ȫ@Dv��"m�o�:���&B�ØQ�K��lZ\��^m(�3ݶs��������4�
e3�fB5����˚ 7y����lƌ�;�����o��.zHa0�\�	׬-&4����5�H��u�u���oS�P� �gr���0�יUU�F��
���0�����+9�r��M���=�}�Bb�o��m�;���w/��.���Z��ٷ@�rS����ҹ�`J���V�3�G���@��� wR,�hp�b�,��X�Hu@���k�x�gz>��U��5u=���c94�^�3�&uw��Q��[�����`y}�cV�0B}ڦ��
bX�s���v�$;H0�+����U�J�}�����Z�L�������&���k�Nٖ����V��ٌj	-���]E"y�C譈	U�&��\��{��{�삷r5���C�/���o5,f�ƅU����x,�b%�����[�i������f`��9�P!R���CMkH����*o�{����CEҌO3�p�.d��B��q4�P��OlAlif��#���8�C��3����Ĭ8��ό��L۩�ս��J���Vʭ�y^�ʭ�%e���Խ��>�m��NUU�ń4i(R��q(�,¤�8���qdD�F@R)4'�:�[4��(>ߑ�h�ash�p����VQ��q�j�1��<5�Hd�L�i�!lAf�MjJ)�&Г��cy����O+-�☳�̗���QHU��¢�E��M��[(�}�J���֓���ӃB���:���WO2h���d�%u�4�!��#�#Ư)��c�Oxpܸ�c^6�Q� Ju���>��%JӾ����'r�k��Z�Q���4�����mB�F�_[���&j�5��
��|�we��C���:�4��R��9�V�`c��t��"#����4�4�\�j7����p�����_;�W��I
����������i���N!�ڪ�芤|�!��������i��o�+0&_X?�2h�����hO��
���`a�E1
�	�/�JO&���v�t��*��$K�^���r����X�J�>
�dAXq2���È����(*�'ʪ�- M��镼2�y����eڪ]F�\��*/�ou�T*K��1��w&Mg�#kҒ
E���H���D��,wRKAaiۣ�Zs�Rx�7�w�o���>3�^y�v��r��܏���d��N��J�[)���J(�b��V�'c�����n�͞6��--i�D�<Zd"t9���m�]Пf	l}�z)����m4Rn�d�~������둾F�4�fB��g|�1�w.����qKsy��'hȞ���x�X�.'�7���~r1Ψr�c��d���h�k��}{�����R�D��"g�s��S+��w92	��"�lei�K��>Ab@�㳌�w��ZOhu�L5�>l�i$E�|M���"Ff���޹m&s������j ����6�����>;Z���Vol{����G5���_�e������-�Qx���᥃e�0հ�T�H!�-J$���'�}Йy����G.��p\.�9 :0�#�#���X�#��u��v�y��Sl4�^��&�V�$Y�2[Qڻ�@X����wy�~�fYT�xAnL�p�����	$��_I���^6�P.���*�kp9�x�OnCv[D/v�0.��cîo?��F8֤%�Wu��֭�d���{|�(�]�e?ni}������Q�)@i��V��0A�pŌ5���Მg������-�P"�<btt9����Z�~���I�!e��� <ڳ��1HV;�ho�|#��j�W� =�\�ݖ�9+9W�UQ��O�W�!�����=�c��!�W����3�3�������c?BN����rHzV��yY�u�n-�|d�����^�
�4�#�h�'H�y�$�
I�:���11Ϯ:��eē�tV��Uc5��c�a��C�����_�g���-�e�f�aL�k/�������܇�?��T�TT�o>��m������L��Rݍ	��N�����zB����A�
*�U�Wn�������뼬��EA�/V͌��As���e}hD�+:p�6�|��K-���Nؐ\�kwv���}�^un�q'jZY����N��[��b��Y����&��p�{
4�k!�l�m�z��p�(�j�)ncS�l���N���L]�U�.Z�2]x�w;��w�n��-c}��j��-��[�!��s_bӪ�5�՗`�}���t�cE�D<��P+�Vͻ���WL!���f<8�KiI7�]˵q8�Nȵe���]�r��鷐Ki_���|�`ۖh�b�RS�쩻k<w>�ޯ5��C+K�)/u�̆ՙ�Sil$�d�.��%��«�+4)+#
 R�6�QEQ$�qBu���[�m�?w�������hDMDDDD�"nj"nn""" ,��Y�&D������؜� w��m�e����������ɐ�����Y��09m }=�z����K9������52d�DDD�=����ww4�	�D��H��qH��I�d���"� �0SI�LE�b�(�q��QE��D�,��&� 6�n(�����[�$���0�F�8����(E�Ʒ�6�Q«�y����Hh�3�2!I"�8l����Տ�����	���m���y�g���1?4���(�U �(����	4�oɢѯ�~�K����iar(X_T��)�Q6J��!���nKx�a2��"�����ʦ�Z�["�J�u�˺^S΂� "��Jڮ5۲)Z�;IX��˺��J�M��R��.��nհ�&�y|�P�M�����M�	��į��c�/ZӶ+W{�ҹl������.��-u-5�-m<���{q>�pN��6��[��:0�c,k��٦��3�#��F屔ἂ;z���a	%��k�ۆ��<�W���	��lPaf�36�QJ���iP7��.˛�o�n���{�B,��3�b�(�?$�J�a�J[K�#���Ŧ�a#+e�9�{ne̘:j�X{��r�:��ӆ.]����3��O'Wn�M��)7A2[��<g�,�|��aJڀ�Q�DJ-T�*4t� V�ba��H�A$8�ֵW}�Y@HE5ۧ-]k��NL=֭m.(� �'j�]�]0��X��h��w���7K{+�͠{M몰ʐ(-���>�7if��B�JAm&Pr�/j��Pi�.!(t}Vu*�4t�
��t0Rְ�����Y2�ʭ�i�1��3;zh�`��m�YD�UcqTB�Ǒ(CYc���0�q\MQ9���ZHg()[�r��̚j���0��K��\6Pj�ݣA�-W0��h>�ω�ά�Du���!�r�m�c���E�Eۡ2��W���	P<:��0�q�ú�-.�ҩ^�&}�_I�dh6h���Po �['��]#���[I���١HT�c�D��3��W�u<������娧���ӯ5�-�hd�ݖᗝ�y��o< }	�"H'��R,�	��U5F#�_M��ĒN�5��ݭ��{G�δ:1�繬k�����U�}?r�xx�~�|׋eI��m��ǯVu�k�=�8�ϒ�u�f�v������C�$�<!����| ��u����Y�/Դ��������f�"�멋���i��!L�]U�*"�,�#��&�k��o��Uk�1gL	�P5&�#CMj��U�`ib��>]Y��FR�O3� ��+�0��2����]�����Ӭ��$�w�n�������]n�B&Ù�!e�[�ɒ�<۩=��� �>ܪ�REkV�@{h�3���J�M�������1�tzoޗ	�j���t�L�MW�E]���"�+�K�X���g6����V2.�ō�#�H�jӉ�M�e8��+n��fD��Ai��(��2��a(���E\Z�K#wE��}A�V�QruB��y7]���&�m�L8EJ@7��ki��c|�:��m�_;��2k"6�<~��E�`w���ba � ����v���J�^����c	Q2C�O޽��p���3���#�qn}��J�r@�˯c�*>����/9C��5��L�Aֈ:k��Y�X�rLk���*�nY�`|��SBL�l?TT��M��.�n�7��� N��7.�a�1%���P��1����N����ײ}��P���7�xH�b������ZģC�Ǧ#�iGxQۻuǀ��˵f�����s��b�~B1B=	�n�[2V�S���z�t](e�9)Ah�Mf��h�<ꞎ@�]z��)�;-+-#��ޫ�S7�g|�.���E۸��ݐ������hh�EV5ۼlڊ
�I!�"nZ۱D��Ǯ�%�L�h�'nuCc#)���\&��h�z)�ު�}�#�([KƯZ)�Y���ja����@L���@��h�P%krH�_�q�fz�ƊجN}��C��| �j����T�Z0��ګG)��#�}��o���seo�4ږ@yw�3��)�l�8z����Z�6W�fa��F��K�O�l�����h^�.'��g�No-ǕH��so&=p�!w�3s�۝��9Q�)Z��l�=��=�g��6������襶M?�>��h��2O��$���U���C����홊�r�����i�x;�7�b_+��4\DV�Q%Ҵ�P�)����A<�mv}d!����!���nE<��W��}��v|����Ͻ������<&��w9���F�!��E�svњ�xx	����ڏl��L��h�J4�wz�.�w��$s�"S(`w���ʃ���ݻzWm�F���n�v>�굀O���![���j�� Ir��tN�g��@��*u
>>1&�!{3dY�����<tt��]�M�Ն�:ZD�ep��z;`�n�܅Jl�Eʈ��0!�ϥp��tw3s#�&ny9�g��1j�1:�f���栌
m�mmj9,�1�=�ђ*ۀ�і�������
"�����_��R��pshV�B�U<���?xJ}�q\$l*��Q馶=Z�%�?��5��'3��>�/�	~�s�%�֢�f[+�l��
��̕����w��Z��>mR�[��A�{��r��7�ڑ#C�=[>����p�ͺ�U �V��d�����W]5_Ϸn�h�U�a=a��v&D����KY���b�f����B��	����c;Fb�-�y���k�t[���yGw끾��d��3�2�����Kp�{Dx�|A$=�ɬ�{�y�R�d���ǩ�;k)d�g��;�se�E���y
9&�-�����h��=Ӻ
o�LJ���}��{������c������d�N�wP����$�hF�_�<���*s#]҈^͍6`Lځ��x;n!vJ%+D4��-�_ҫ�w� �ņ���v}�����;Mm��'���y�׃q�)�ϥ=և� ��s-��̬�C6I�1<���dKw��(��N:��F��Z��zԑVՉ�=�p�\�.�};w��%�ǔ"���e�i��΀�i��5k%ӵ�xϾњ�k��[ͥl��~���=�l��^�w�;���96gٹ���q�8,�(뻾T)�s�J�ͤ����X���O7)y'q�A��m2�1��M��($!��ܬ5�G����
�x>�s�҅2�e���'ka�5{�L-����=�n���;�Yl�C����\I5��ƕ��*�ii2q��g�*�m���)��z��26�D�_1I�l�<��Y,A2'S�G���i�lb��UT�+�m�M�����jQK&r�}�{dQ�A1n����BL�g Fu��H�nn*�L�|U��._��p%�N�� ;Z�mnW5�۲
{(LJ�U�8xK�]�A�N�[�3�N��P/�;�H��	Ͳ�9LD5j�^��V`L��|O0^��z:7;�m�		�I$9u�D0fK@�l���n��K!e)AVZyك�"ܶ�B�Q����30�,�ӗrY��HM[.��Z�OZB���WhX�n��8�l��Gv��X�r��6���PRWS쾲���3A�/�����Y�\ǋi�}��k���R&��'F�"s-�*ϋ4���1�ۻޞ�gu>�#��R'����byuUpn�wZ��m��MWƽ��JoB��)��l;c�����^K�C��xx6��E �(�Q'Ľ4�b�"�̼h��i��c�;jФ�zOI��
x�Y���p�	��!�ϱ�vsl&Y(>lƃ����9���x��m��,�4�'C�+�yu���
��\v�.v`���=�F�HBֺDj�C��{�g���y���l���9��dV���,B�����]��D�!�W��i�hu��� �0��k��6%nBS�r�Ɍl�*#5C����2/0�DTa�=ϊsu����`�E�ϳ��IE��fD �%q��w�$����Zv�P)�`.� s��F����8Y��ڗ:W���$m�DM�5�Mk01�*���u���1�~�\e4x���y̌�i�(YV�0��"B"m|>������돎V1����z�Wn�Z��qy�(��DT����3�X-r�̉�m�uhT��$�X�b�Ɖ��50�@�e�n���(��o�yo�&�(XL��nlB�)Ac�-��^z��pђ��@q$�Q����D���Ǽ��۝��[�$Md)�$b��mX$&^�xTЉdَ�=���jУ���Bg�hx	��(]A�"��J�^����#�?r��[��*>ܤȻ$��;���wx]�15���DI���ٶ]����7{��P2�A?S�{>˩��V�yq�h��a
0#Z�r��!>���p6r�;�#��e)�	SU>�AԂ�N����'=��������hw�UK�"�� �;b��7��q/.iz����4����A�r�I��G;�R
]��(�DEC��.�r�)�� �l^ɽR$�{k}S�WR�U,�*@Y�Y;��k��/~�|��nn��e�m>�������짅����8��*V��+���Uڳ���!�����AeZ�$qy�!  �2kB�?
�ɏ&���{�����c[�s�q��Ǌ> +��vS�����Q( �p����L #l�v�tu�m�<�^���,ZZ�4���"Bh]��H*E����\i��}8"H��R�	ب��o֠��q��h��W�F��41�1"�޵���Qf�)�����oѹ�H�vT�]a"e��X���x0���}݊e�1g?w}���4��D/L�3B$!����˙�b<*n�~���7�2�w7�n�}�t}$֢��&FKiA�$�u䭲J�K��l�E�=�G��b�\����0��p��m�A��@��1T��k��sdH��{ȏYx���{��u"�1I͵�!W��t���+���=�@$�}8:z��������{��}v�{<�/v��`���4FZrR"i�ڂD�����m���n&�i�I24�F8Qm�؍���P�VE�����O�#�l��e�5� �@�Ȥ��䩯K!0BI"�%=��l�ˮ�!��u*�5[YbX�pJ��9{��f`h�b̰�8P���� cr��JdRx(��\t;��@��N�y�"�z���<|r��
�M��&�����.�n�2�\�H�mk���x�gЅJs�M�
:��:"�׌�ê�dM0�ݱ�lg�te��3�86_`�G4kY�� �hi$���+k;��uo��0�Q>Ke�I+T� �I��!�Ӧ������T@���Jc�3|"a�A���{ꬖ�p�td8�s.�O_�}-۱L�"�w�P�RgtXE�ᜬ�{���y��!��F	A�L}d!)U<��ɳ�F��Q��m-=[={�`�=��!�H]�������8�fZw���*!f�����<ȿf}3s\�W�׆k��=d��;hʥ�kk"RC1)@�x����.hy�j#B�#i*�ō�x�&P�LtgQ�f��{�0h�ۜ��$$4�JgX�`��)��i&��C����E�g+x樽���-S�q	��P�����hf�D�U�ָ}Q���7;,���]�p�	ӗ�o7��t�MU��/�0}��XIv�w~�<�ػ��/�Xækf���lc���NW:�`�6��,��X��g:���mK�,ΠCul�kz�b�EZ��p��hB�G�ڌ8˗�Y�^<�[��2v$pU��em]1On�+Ed=����w��2��J�4��n��̆�#�|�:��:0Լ�s3�����UMA�#��g���5��N�㪆��n�.�t�9�N=k���5���n+u�U��g�+6���M��J:��=�Eԭ���o��%�1W�or�thcJ�bϼ:v��ެ��!j�7�q�B��:,$�у=���w&�I$�og�l���vvvYb"[}_M�[ ����n�րԍ�{ܞ���̲�%���������y�q�Ae�������7�3   9{k��D#���3��k[�jj6�����_&B$:�
 %�LB�$"PE4bP�#J9	�5)�<LLׄ��b-��DJL8�		��C��u��~���e���GdA!E��+�4���s�#n6�I:�=O�l[�$��R�&ͭ�kHc�|�,ԉ�#�S7S�c��\+1������P7�hQ7w$f-��jX,_BOɓ�T���N޲��v�iY��2�Ӝuu��EKy�<ּ�=|������h��Z�;�RxÙ��s�}V��F�����Z"�Hq��}2�UƸ\X9�f�"�i^!�@�K��U+�E��iK���K�*C�v��s��i��vy'}�<��Va�/U�C�B��yR��\�����Y݆��7���uU᭎�+����/"�)ص�Qj��W�[5WN�5�`zbw����4�[�xƂ�C&�ß�.�BI}8P�q�룎��G��V�fUk����ʃ�9��[�τ�`��s�.ʫ�CRa=Ĺb3��d�/uYʞ��s��n�*�|%ܾ⒬=�ݘ$m�6�G�}��� jDct�!�)�|%����-҉�	y�*m?$��a��_J�4Egl����9[�$OS���z�gbdjo#�do%mD:�K�lY��Fnر=x|k�d}&�t`�$��S^��{��cݏMy���o6J6p,FC��*�o�ŋX����ӂ�jJ̴�V+���(csR�����	ēI@��I�ƪ��\xDqK�YH$e�#HaD�6w�����p#R��a>@I�	�h1�}BȏJwjh4Bh�F�|ۆ�X h�[��hG5�&�|��ڴܻ�U�@L��yH{s�J!Uu�N^�w�rZ-0�۱���a��G��c��,��J�B�A����-�N�c\'V;@���Z	�_�V�r݃�b4U�ѕA����֞u���$�%�R�`�����{2�O�k�5�*���o[�M�ۄ��N���	bx�͋�RM2˄��hm�E��b�S�f�ot�&�;\BSN�+6Ҵ��%)���rr(�:�Re"QE4	z�	Dz㓫e�ýb#���;PѴ��*�Ë3�M| ��q��x�6�T��4�Pad�:��k4]Bҷ���۽���=�nA��@��1T��"��T�{"��xε�W�����,�%��@��v��=�+�ೢ��jw�UHt�E�
��ˠ�c�{t;�DFc����MЗ�+O��t�I�BmN�a(-���j���	#I!���
������g�ǂ��?xg�n>M�Δ�fC�P�����2`:�f@��0}G=�RE�a���/N�ۿuT�K�n7��5�0� �hi$� ,�|��{̺���"xU��e�T1{/	C�H3/��3v���;���˘�6��v��F��m��VX6C�ֶdn�Dfie)��!ʿ�����D�3���7�{�&�軎����☌to�f��a�)�woq ��n�w��K�	�RD$UH�~���|HM�$!I>�b% C("v�R��lg�0+s[1��0̜΢dD��޽��"��ռU
��}��L�"�Qƀ�J;�=���@��#C�fhaRB
!��{]�\��Gxy�3����%��'�|F]iqf�WSÄY�<0q�g��3�G9���څ�o���tY��E�ٟ��}�3���	0��9��a��S����]R�D�=����o��8����2����>���*�}�i)t��n���y���Ϋ��*��D%��\5���-Ѓ聍���	��Mj�>��宓 ��5	BP�ɦGxhsٹy��Mً���S+�DT��K�Rt	@���X�y���k�Q��n��yP#�����rD���s�J����y���xۺ�c�~Ư��Ԑ�iд��ILo���k��5Ӧ����	�A*J���P����w���.�Ϫ}�Y�ZG����2��p�g ��.v�v��y2j,w��Z�!m�����R�H ��(��	/ U��	�b�j��o��.�A��i��f�i���CSA�P�B(�I�	E�����a��fK����/:���m���\c�E�)$J���t�* G �0B����Ӛ���.�_Y1��0̠΢dD�����X��{ZHrR`��:uEAw��C��QDV��@g��I[�'��֮���b�&kB����Z�e����o!��5�[9�n��V�h6g�d*4D�����.*ŊM]6#����m25��ta��QC�=�A��?�#�� B���f����PnCШZ�C��\=������6��4C�-���2�+a�iT�,�}��MW"���!���EJ�$��[� �gd\ח:m���q	�ձ��yf�YIE�27�� C��Oz��U.wb�3a.D�4���n0C�7��bH�!&!�&�)�e0������'E��<���Ulޕ�(��e�RW��eK倲�#��4|�,�USCl�!i1Y�hX��8�B�GKxm�����h��"Cu��
ք>������u�%�K,���&�w�9���i�B{��(cd�"��2ڪ<a�x2]*����n�֔�&��j�W���S$p�"j6��T��\5k���|/0b"��5�0�=뱰%H��Z�	!�
�ȆC)<��-ָ �rm�Y�A�%qQ΃�!�\����QlyI�y�n�r;�F�l3("mJ1.$b��a�Ө� !�Tw�e�}�����Z����I�	��f�𱆔ssߎ����n��(w����o!�m��w�ؽ��
H�
"Ah]ǆ�6��|�£DI�R�H��sr!>��"f湙�+�
�}�5�%ii�)���-fEPl���	���
wS�}7E�Եz��4Ug���we8NDڒ6l^��C2o7wd$���r�9�f[~y1�K�.��Va�sY���>�F�ʔ��uY�-����-J �8p��D�H�	b��)-)H�IwR�y����:M���=�8w��j?�����h�DYP`b�� �c	 B�y�����מ״��]bs���,���bI*�����f��a��:��Ԫ��"� 0]���ow�
!-�;"b4'�A��k�R}[��M��ɰ�q�M�"�_a(s\���C�^9�Uϩ�A�Q�6V�NQ���	�.� zi�� �������SmR���N�X[���-ϨX��F�����!(?oK��3�C�O[��"H
����yA�[-P7[�����A�e8[N1R�E��n�b���ɏ��o�\�[Q�֜Tk2�"�E�kQ�`����ݯ���Y�{Q���}���-t�4�/���w&��*x�	��<���%u�
�<~��)�{3����ټ.�� a-�����}�/�H�ͮ�o�� 6 n^�\�u!�|v�:Xz*�;��J��fXi�AwV��K�Ra��2$2ۆ�c�JB�l6�2(-��`"����i��9_�/%A�D�1
�T9�C��� ��yM�.=�̲Ii>c��m>"�V�FGB�q=��<��FA+זR�	��!�a�\;Xd{�SS�۝�|������1+XI��S��ް�Q�~�:�Auk5��z�k�ч�k�+/�}�D더c �،~2	�������C���W����(��	p?����O?T��dyY��r�f����JjϨ��&�z�;�O��l�n�aT��m�R�N�Ff|�����x�Ӯ�>�x!ň�fC&�D 3���]�K���D.;�`)r���l���2%��H�c��X�{��A�qd� ���5�V�_7��q�])SPW:����a�f�J �A�	��ȼ�r�CSI�\���R-����_k��v!�%���u�ڽ��ǓhP>�!�<��a��xō[p��fX^(�
dHa%!����j��-��[.��ǐ�b�j�A�jWC�X�|���1q�!���+������^��h�* @\�,�}�L3'#|1Mʱ�j�
��E��a�����QU���w+bI��T6ou���D/F�����xG�����X�\K[�r_��1�y�ӟ1ۆ٦���`џ%���/�ka����Rլ��	`r�sڂ&���#Gd!�����1cw?6!>cn���!d>�&����]�Bm�"���BAU��F�*��@�ӯ,�<<2#S��1��~�4��b
!+B\���B�I�{ �$D<2��4�Z�2M�P�`G.n�v5~��+7%��7��m+���7Px��|���0Ƚk$��������fea��U{���]ũ$w�L4h%����\I�d��i(�J3+��Yh�VyĄA�FH�%	*$	{܊cz�t�n��x��on��;�݀ �x��H��g�pa�m�!J�["�K�,�UT2�5u ��2�-	I)�۽�޷x��6W���H�VY�p"*g���%T."�J�Ag�==쀃<0U����*����n}��;��O� ��$�-�U�I��ϛ�E�����i����׵m���=DC+�6%�S����N:$�Qr��y�m��k�\���;d���g���eN�-��,�ǟ@��+C��P�}-��L�"�Qƀ�J8r.m�Q��=DY��AWj�2(b���{�*��R#�lBK&�͖�:�z�h�z��Y
�$p��t+=�)��J�L=[�R#��i����A��n���8�(�ş"�L�y���@��1MM�#6X�������ݖR���h����߱��FU=�Kv�%4n�r��oI[E�ӷy�}��E�U>��1�<��v����z4hKD"�y���L�R'�u�Yg	���h'�i�K�m�ŃXr�d��c*-��:���.��Qq�g|ќ���j���H5B�IL@�%$XAQ�I6��A
@] Z�I�yȋoJg[���S�� ��\~�D+P���b�� �g��g\d�i�^�4��D%qF2�LG��1�@��+���u7C���+�5�d��x@�Yé T��^A�]�`e��m<h"�ݧ��P�>!�ܝ7�q�I4gwwFw�3��6ၢ-;)�I��h<=���G� ��pJ,���c�c�#)o�m�X���Ӿ�A�)@/Ւ�$�$�Op�F��D�x͐�
&p�f)��9�V��ɏ��X�R������ڔbV$=��O!A�^L��ʆ�I�u=�H�/�.!G��Na��g}�#�|�YJUO���ѝ�H��T�����[��=����-��z���p�N���>k������w�
�d2��6n�����#a,|�d�O�m�]Mf4ݷZ.�E��Q������?/��Q}P��5�{��]�L4�0�2SOP2�uAId)l&s��|�[-��R2v�����
�-�HD�-q9.k/��^#uY�J�I�$����ye�rEJw�6<6B�ӱ" �L}SB�g���m�٬~���o9�(x.��kQ� ��0�C룔�fإ��,��۽�š���)��(��;�ҊC�0��;��=��N�D%3�6�A�@�xe'� s?hK�A� C����{���[L��us"\m/�����zD�عE<�.�m�:P��z�P$9a!�Y�gO�/{g�ۼ�	t����7J0�R奩��3KOxM��g�\m�����C!��P|��]�/=�g�ނ�7AU�d�����n� !]i�٘�^^Y�s�܆��/�Nz��z�)c��ר���ƴ�2�x|�U�a)�ZM�����ښw;�K-=��1Y�זL�ئ�(,aeXf���SZƨsV�4��B�CF�u�Q2j�ʓu�&�n�k�m�(c��9u��w�e����o2q�K��%�+��#��^��ʔ߻�Uor��;&�NE� ,-wC��^��ꉊ2�vt���F���&b�sM��-�����E��߻��b�t`�\�؇-/�JrBo�#5�k5���CfV��F�!>Ϭ=�R���O�b��c���HV���[c�q7�Y��U�<�3�ɳ�j���D��4��[������F>����>'3�C����S!U�>i��oh&��h�ѓժ�`�ʈ��E)T�2���F}�p�����t��e-y�wsv}U�整�d�f�d�)�LCm)�5����x���
�6��9W�/U���B��u�{'*i#� �a�FR5S)�0_uT��A�Y��8vLĀ���<A�Gݵ8�}�V���
�?^O�+C��3c�X1�Rֺm���/�[��ư�%V�t�a��u�ӕ���1�BJ&Љ$��(�I�O7�{v��C�w������Q��DDDDH����������e�v�2dȖ�������-�����h�s��S��`~�w&C{��ԳZ��2�CP���� ��Ȗs1��ɫ%:dɃ0`9��j�sZ��U�
���L ��T�Q1hqr�IB?#�d�1�m$j(�&(���Y�0�nB�L�'�a�цH�.DL�&�l�HEȡLD甍#$L1�aη�s�U�n&V�j�\�w�ت�݂�LB����M���"l�Wq����M9"-�*�Gu��c�T�{��M!��$I2�iWJ���)Y���n9E��Q�)���'aҨ\q2I5R)���fDa!0�9��, -E!��p���=*S| �ԭNV�6��=�&�g�`��w�+戶�r��/��L��H����;}�s.	�'p��NnG�51��to�iLZgy��i���	Ș�p=隨k{&�ڻV�λ\{���7��gSٳF�/�87wo&��.�wo�x�uY;�����`1]T����y	-6��#1���r�9V����7��*M���5k6�T��bS�:��UF\����K�ru�1����u;�<c!7$&W^K��z���{y_��㲝:#l֌�>�Q�f,����2�۝���/6o9]8,敷6P��E�`X����c1�n�E�M$��p��K���`H<��҆a�Ԧ��W/%r��C5U�1-Q�G9�����#A��,Չ �.��6���`Tb�M��Z�R%�a�0[���{��n���Į������$�F4�AH>ΚB��h����پ��������90d�W�f8�CEJ醱�����d:���6���`�!��� ��j�ڰҘ��9b!�U��f�x.;+Ic��r	ońUF����xV"�8����5t9Ѽu�)�]�ľA�S���]�\ �#C��ޫPSJ�\Inn��ls[�A�O1 ͅǵ
5�s+�aM�	v�՚M�ٔ���*����1���5w� 'e�m��V�I@NN�� ��+6]#	��j;�٪��3K�dل]���5�ywQ�39�|�r�18M���ez�� v-u�땷n�﷝oXƻ[�xXi�
@�.�Y�0�� ��`L��I0���Ȱ��sTCNsT�;��y�π�9�2'"h'� �;$+�a;��������:$6��м��y�3G $Q���6HB�ܦ��^�C�r��|Gxn�03��$I�q^��.�r�8׊�i2D�(98�,��'i8��$�^rS$w�۩�ר�@Խ����عrU��-��=��T�����T�UP��]�96Pv�@�V�{$�/h��R��)E!Z�T�������Q8�&�8ЮPs遭��'�u�B}d��,8�s���ӈk�\e/bC-������G{�o_ߥE��^}4R�^&,Gͱ׬D )�Ӣq�Wsf�W����@J�5&�1tV	sp)���|�'��lP��������s{wy�!K�=m���`���(Z�	q�iI&;U{p�Y9ԁ4�FB@n3BH�L8��ē��˥G �;;o,R�v�dk�%��oTt|��0�0�W��r"�d��q	r.��S����ɲ}4a	�A"P��x���w/�KiX<Ay0�:+.[<�X�`�q���}I2�$�q&�G���đ$B;�0�Q(dKu�I+{�f�m�޹�=ᙺ�I�!ōYj��IL}o����ޤu�;&VGZ/ ǥBө�>�}ږ< ��W���E'4��D/L�a�340�!�ˮ�.gы1��ڡ��LD�\��7~�����{�͎��_;G�d�	�����߰�0�m���=+���.\=�9À�l�+XIlԱ�G��cS�4<�Iu%lЙ�-;`�a��7�=j�������� ���߹��b'��)�g�HQ	]H�������u��ޓ�ʠKlGD�~nf�N9�TIB��y�%��l�N��w��������2���5!j�u��BB�f�.�1�.FӅ��f������i�)�d�,T�,�Io��Vn�5Mn#}�7\�:��mL��TYY�Cp#���XK�/x�kO�7P��CU5X�&���Q<���ۊ٘F'��u|��L��H |O�����GȨ��RU��;�J�yUhSb��|����+e�1�6��`L��}e�t���l6����r
�U'AN�=pi��HЩX�Ĺa��ِ���ۆ���{�=Z�CF�<�t�aFD���I�Kȩ���x{
�|���yA�[-@/u����I"��f�IP��uI�yd��g_��ew�o}U�,F�5d��-$^g��~�-��_�����(�JC0l�w���!�S�E�0Qj���BR�|v��o��̒[,����D��S����k�vS/�_�ܾ�`$4��#��CJn� 'Q뇰��L�f�K��g|iݟ������^�1��U���4A��#6��ՕD�>��Ć�}vZ�]b@�IdA-���8'"}��/n�t�EJ��_^ڒ�T�z��,�ksr�����IM&YH)]�����!N��fj�YT��F��5s-#�P��C	Hk�i����@�4ɷz�I$�ʢ�n4�[�(��A`��P�]�2�mZ�a9h����'��ŷlA���5h���.�w�ȱ{b�3��cˣ4�fإaЎA���a����
�x��t�x�G����HQ	m	P9���~���VGt���P�xe��W<�}d�M�1�Y ��j�\����!�c�(@�R�oTk��6f��>����UtQ�ŮRD�q��(�b~����H��!a�@���@�*^�}��W�K{��m4ְ�"Qgh$� ,o"| qy�[�<z-M��mz���B2�D+�a�W�k]M���()��,}��L&ND�O@��O5�5�1Α�?��25�� ��'=(�S����DȵՓ]��5=�	�
k��>��y�x�2�6i*�S�b[rF@����C�����G\���ܱ9U���W8h��6L�y\a�:�S�v)>�ݻ�����>dSC�Q��$��MD�6|�"n��F"��2!yœ)m!�kE��D�5�PT8;�8J%j��9����~F��e¼C�:�N�����#�0ksWQ:=�g4���a&<�:�2��P�4�W%����z��V�P7/a9��9q�.[�2{s����0����; s��@+��F�n@��)��������'��9�~ė.��:!ht#r0};�] α��ڄмdE�,�7w(��T�RhW(9����f����Mh_��<��Ɉ���Y�i ��^oq�1�6<a��J:�Bwi�B�@��*�N�㹐c���Ƕ
�2���<���{�P�B(���(ДY�	!��~�a�����{��.me-�i|XӹA�Ş�*�C�o��|�1.��֕�M7�z�T��"{K��%�+f9Y�zh�F���Alj3<�0B�q�㻝=a�U$$9�!?���m#lƤ��k"�QFM 8z�6�c\����%�rq��lh'1�
�̅��P�Q%���,��8[��T$�/��r��lÌ��8�m�8C�-�n��{�I�ζ�\���{ھ�aq��Y"-�c���V@����T����j��]�9��f�~E�Q�&("t'� j��A�p"JE�3D�'7�>����ƈ#5Y�A�UHYxGʭn�3Eg�\0���=���A�#��W[9�m�<D�0�J�In��a;�;���v��U�χ"xv�PA/`���9q� Ya�l82#��w^�O��Mv��^�ʹ�25�Ӱ&�*��S��������A�����0�A�6���>���=���5T��(��L����a0�L}07����$�8Ȑ�8���G/?V��d_�b�˪���ću�o�؍=�w���n�N-HS��5��h���i���8lW�[�Z{C��>���V��fJ'2�{�ٹB�D�|���O�eH�h��<s�k�b"�!6 �f�ل���J��T�j���na�{_�x����o2�ZX$��-z8�>� �����L�D�	��A>�E�A������:+�|��gA�?��I�$a��v[!�<�����=��WZ����!6�$�ѨZְ�xCB�l	PG���I@V8��2����g���n�͂
��PřI"�����I|�E�y�n�FGr�F�s}�h�0����U����ر���>�z�b�RV�w����%��G�^��5�!x�հ�z=�̮Ii 6dlM���6�,�������!��+��A*u&eXrof%��&"��Dw�h��q�$t[��)���|M+#L0r�X��.��c|��u�2 ��͈%��(���M�lR��F���
p�c�p�.Jb�̣4�r��\�����5j����r��T{��(����'�i�b���p�c�T��U��ԓ��WT.Wf��i�V�����{η�[4Ya�$'(y$@�Q(D� ϙ�h����%��-o^����N*�gZ�F)
�;�]L6�^�.}(��{>�y���C�|�|�v1|�����/�v<�~<����Ҽ6[k�~�J��<'�Mxk�{�n��;�\�5B�XH|vd:m�B�������\�M9�d9kJa���Ϭ2ãy���*�7PJYy3�^��p�H����t�P}�{0�F��<ޙ%T1
Z8�w��]t���n� P\��G�w+�]{qoִ\�#N����
X���P����ǝ�т�f��;��������Lܺ�l�O�sy4���1N
�Vu�[9rnGDҟ����;����+$������1� @�!3�;]ת�v�1���}�	��:���\sm��1W}��&�.�1wS]׼���k�p�U�'s����Z�x�<����چV��η����H���� g/8d�TA`�5SW��m5���p����/��b���lK�0�������.�)������0D��Z�a �h�4x{�1�{����r��EBF�9�
����;����ՔY"IG�&1��8P��8�N�b���ܢ�R mH~���D۳�6e��w;v�A�9�@רc'�m��b�M�����Y�j"g0�^:���G�=:���t#v�8 �Ԭ}�8�!�
�̅ΰ�@gm�x����n�"Ȧ���/*��ZdȔY�	#�����[;D�&��W������pT���;��_ $t�&�j�H�Ҥ�<?��f�3ЌJ�Rk�u�=-���H臊�۸'��wR��T/�ςg���l#n���Jʵ�㌲m �^oYB�<��ץ�� c~�m���T�]݋,=���R1q7Pȋ%8"l�:����j4�6�D��I�Ȥ�8ڛڊS9C�a����jMޫs�ߊ����GÈ'�I1H�PsДs\�BE�Q��44�[C��{�Ёj_UѤ���v2cA ���݃tnaA%�a�ٽ�
�$�T�"	�jS�%*��^������ �f�#z�r���n>� >�lK�dE�0yH%���x	|9[��=�{��/����A�z&�#�=7U[k��Y�	�aau�&"_A�Gې ����s,VCE��t��L�y���
����5��[Gxw���e����^��Aܢ�SR>�˽����Xw|�ĕ|�Lb�Y������~��3���{�|�8��E5��q�kɼ���������czѳ��Ë0R�Q��!��L"�w@]�b
H$������������T! ��r ��!O��c"H�	$��Ba �%$���!I Dd *��P	
��B
@�d�]�HAI$��������I%�BBO�`$	� ��	$!H� B �$9��o&�*����O�$ I!� �Mq�����_�N?˘����N?�R����v�?L��O���O����P�2 �#��?���,��������p$ &@  ��Y�~����j_�
C�������~����?���7��'��$ ?�������>������������~���K'�
����C9�LCt����������_��~���_�?D���� �W$!I E)!$ �@P! ,��$#�Ā� �@c c R�@H� �2D�� �#$A $H	H� � � R�d� D��@
 �2 � P$��$B�
"BD�d ��)@A�$��I	�����!R b@d@ $�$��� $�H@� �$ �	� � d@)��H�D�ȐI	"A�$ �FD �B	B$�H2dHB$�$$ �H��A"A� �0�A ��@�DI$�@��a"A!��A ���HA�"H0�FE ��	H)	�@`2$�d@@H0` $@@H 0���(B0@�`B0@�0Ȑ�@�D� H�b � 	 	�?�I(��@d$�AI��$"A ���� $BA � H0�#$H$Hd(���A P��I �$�`���d`2A� ����$2�
AH �F$�� ���A@X
AH
H, �"
A��(E � ���d�$L�$��A �$	�A�H2!	 � �@"A�$ � A�H I	$���  !	@H$�	�BF	�� $@@H$H�@� ���H$�@a$`0��� �H20�	A ��DD��A#"D�	��	� ��bA��B0"A  0� �H	� H2@�A�` 0$H$H�`D�#�d	"A"A�"D�D� 0` �D�	D��A��Ȑd�D"A �`�@`2 $		�A��$ �$#"H$	"A�d	"A�A �	 �`D�!H H�d 0I� H�� $A ��D	��$H	�� �H$�A�"A dH�d#$ ��$0�A ��Ȑ`��$A� �H$dA �$�Y"��0 �`d	H1 �@D�	�"	$��A��`�`�Y��R����H��
�0 1 ădR�A��H2 !"A�� �" �@�A � @d�$B	 !A��d`$D�	������ ����"�P@P��BE�)$YH��RB��`
Hd�@F Ā�H� � �� ���"�� " � # R  F@ b@c A 1� 
@F �0 "@X b@P���B���1 # X $`�,BH`	���@F Ȑ�!�� 2H�F �$# dH �$ 2�2 ĀĀ�d�HIH��0H
@D��@H��1 1��1 H�`,�1�
D!	�� X$�D R� ,� D�� R� (�@d`�"@F@�1 D�� ��Adc�C�+������������@2 _��!���,������������O՟ݯ����h&? �����?���8���d� 
���J���3.��I�C�������_�Lb~�g�������x�r,C_�������?#��8�G�?�yu�O�~��w�[�~�� ��?W�h�?������~��������@�  ��>'���4jC���$� ~i��h~��x�����0$ ���ș��7��*����Ç ��U�"���+���f����l����O�ka��b� 6�������D*C�(�������$ ?I�����������E��U������?ÿ�A�M����_���������d��l��T��7��@�@��������?O��������~��t! ���/�����W?D����:��y�����1�,�����y����	��,�kA��PtG���_��� ~��X&�)��N�#E���?�������u����������!��������H ?W�a�E����dk���X �~F�1��&'�3����g�~,������C�������b��L��N}8�� � ���@�  nO����>�ΟV�h6e�U],i����X�����ɘ��mBխR�V+�i�m;���W�.�ݍ�k��hړM����)l�l�Po�         :�*�ʫe%Sh$,Tf�5i��m���e4��i��Z�j�-���jU�M�2�MM�hf�3F͊3zn��f�dkV���iVlkZ�����YE���fk[T�V��Q���F��[Zֶ�-��i@[[L��)*Y��Ǿ���d�5l��Դ���ty7Q��{.��P;=��)�M��9���n.f��;N����p��uG�.sf�3J��+X� p��h�֖P�UUZS�*��J�Vy���T�T�O{�ޔ��J���y�P	�� 
�7��� 9��v���� ��fp:i�� N��5�ķ�;�v�$��L�*#R<*�N'8��w7 ��Pv��L�p �cp �� ^��K��
 ���[jI|�C��fԖ����e� �c  � ��8 n��\����L 	f` 6�8 s �ʠ[iE�
7;Mjm��Y�����< ��� �u�� ۛ8 �4� � ]�� >���f� ׷�� k� �t��3�����V��i&� ݴ\ p, }S�{aހ�[�� �w�� ;�� �� � �n t7vj����5��s6�Ym1Jؙ��M�B� M�� ��;@c������& ��x =N{�M�� �!� �W��R��k1B֨!V� �q� �.8 v ���� ` -H� �!�  �ם  2�=p =A:�j>4v�*j�֨SH���T< �a�!��\��� wV v� Z� �n� �!�� �OT�mUUZ�tpa#kj�U��FU[o�� =us�p 9����ˀ��n �;�:9���k�����  �{^���                  
��~��)T= 0 j�����P� �	�����$z���	����
J�L �	���&B*6���i���A)�)��Q�jh3�����Ҫ��g�|���@��Q�(���l��ٶ0��fͰ?�6����Ͱ?טٶV�f��l�s����?�����?���A�+��2���=L�(��/�pp)ʬ���/���Q��r�9B�>�u�$�ѧ��Fy�0�����ճ.��#�\��p����@�5-�t���ȡw�6��d��Z�(v���q4l�q��7zfY���UK&m	I!k�	�:��q#G��|;2��gYeRƂ��,�N:B��n�$�Q�gL<h��@��6z�r��N+��?21�A����$�a��!Vk^X��M�(�=�#Na<���� ��	**:i/Y�W[��3i1''���{l�����`�!ƞ�ѽ�u����r*�r����U&��[�t'vfj�$nU窵�z�-��2%AX.�w�"+t���\�MY޴�iѫ��f켠u)�=�x2<3����^����ʫc]�B�M�{Qi6��Y)�Ou=�u�5F�,�E����-1
�E�ʴ
6iJV��nT���<�E<,����}�|��g<�\��p�46�S��9�]�����X����*�Z�Dk7�V6M]^�ޔ��Y.�:�%v�ӳJ�g�K|D��<�3B��e��������ZF�����Ys./!��3���D+xjS�K�.�[�F�V����2��4���i(辰�鳙ڸ����Ő��ܴ��H�#�{�\XӪ�Yk5&-8���@�8���76Ž�Ψ'lQ���X���
j�����=&�6���Lj���n^RV�v��u�v՗��u
ʠ����fv+dH������V�����+XRN�B����
��wR蘖]�F��I�v����02��&��j�l��57�����-�˥��M�R�ů��RwR�]]^�5!��a�Rx�2%:Ys�b+8z��p�K�pM�EZֆtP@��f̷�ǁ6�TQnbI6��1E	VA�]qEM�O#�2�_&(��NMŧ*��i��к�J��;��=Nª��M�>��<g�93ɜ��gS>[=u����\�ThnGj�����3,�"�1�(�f�x���&�]���\m�yL��BS�-�{�-,oA���)���So�!VY�]�ϒ�W�4�ų\������{t�E�Yi�@��zJ�׍�>�7]��W,�����uf�>��q�Ɏ��Lۏ��6u9�1	4l�2�S�v�˼�*������<�J��9��/\2�:��s�W��Fj�e�珬J�Ĺ��v�_}��-l�k���t�����5���ZwO�l���X)�4��޹e����es�����څڜD�Xv��+���0�c�!�C&^o�����1���UQ��[�J��ݧ5;
~��Rx��X���!��3�!G�#�H����ҢNS���e�ko�}V��� �oev�|�]�8ެN�6��`̈�R�Ö���A�ڼݗ��};�?P�&����aԸ�����(��@� c�b!��L0�1H�*����R�RI5�R*�y�YS"�YamVK�0�7d�L��Pe�o]��ebV��a}L�!����Y'
0�f��z^��$�Ī��ŇMv�d-!3H���i[{s��U�F*�*��X~���Av5��qZ9W���KD��Q�eB�k�w[ �)"qPӖӻ�J��v���U�z�מ�����e�3�g��#��n�Z�׼Me��Ӓ7��bä֚0�/�s]5V�i��fN�eTM�2�H��t��˄��۫6Ÿ�3UH��R�+(�r��%�I��6�د4ۋdR3*��j�]2��eO��>����y�C8����Z�"�i�#�H��b��7zp�L��*��� ��#
q=Ȃ�2ŌPѢ"��OS����z�����U�֦ja���0P��-�fK*au��[<��*��bCR�=�x@�;ϻ:eQ�4��=�Y�O��l��u����n����WUNV�ov"��88��{�iu͸�G/���\n�q�S����u��/e��쩜f3�Ty��s���5ݹb�M���_&�O��o%�-���LmZY8۵�(�akh��Lhӷc��y����%=�h�ei�u.)Z�=Qˢ~Ɩ3M<̼9\GFr]�j�x:MY���˽��_Fq.1��R]�g��l���zضs�j
d��{vT�x (��8afQ��N�<a�wX�%�/���"�6t�㥛6F<I��0�dT��%�,��Fx�͒E�4hÏa�|��V�+�>s��DD�Ѥ��},�]i��\�?�Kxi�Y�}V��a��}S�^�'z�^U��Ӝaš<�o�7egsl�z��JW��/q��Y[��M���!";�퓺J�ڮm��(����m�tgI{.�}2�l���T��Mu\^�h{o��\�P+I
��Q�UE���`���,�fY'�6n��Vv���ʱ/[�p��=��_*�o���Dogs�s+\��=]6�X�#u�����%�S���l��R��ig%s�k�#`��⸴������ڝ�C�Vb�w7���s���={3L����\;���{1'����u�q!X�UqML�b���{x�[�s�Y�/�U���[�j�fKvh�Rb��mb#��*�:r)ӫ�0�BUv��#f"�4p���e�Bo,G�� �$�fܔR�����u,u4��ޣ7���37TVX�WA#g;/q֦�R[1���]8-u�ǱJ��>M	��WU#�.��w�Y���]�yvŞ�3E��	^�W�+��Jꡲ�s0���u�:nn�A-���Ì��
2�ܚ�Z6���3�7�)Ǔ�
H�Y��C9�]��Rom�6�V���sv��N�֝�W�p����MD+]gRkr�� �p��i�� s��(ݛ�[�7��]PBXpe�iG�ݬڴ�V����v���g^�K�7g�`Q�D��S����vv(QN��+睕Bo�S�L���b��dK�:��̃�i�8�����ee@�b�YB�S��̭5U*f�w3D�Re�K����V���<�M�SܲP�+�6�V��� ��3�R�|�ٚo��d��7U�t���+��M������'x�;�x���m}KU��}��I��(�'���ƬX�v1ń�xѪ��$6�Ј�n���f�Q4uF���r���U쳩�jn�UV�W��-j��,��=���e1i	�ӝT��X�ff�cr-b �ynX�n֝J,�m��!��XPm�nV�݊i�UD�B�ڤ����]�FӓH��i�l36��\őZ,aH)���U6 <����d�8��m^uA��]d��B3ם���;9w���c�eT����<f�n�6.���&�����	2R�
���#�����V��LNh��-s��w����\,�m��۽|�9\r�<X�Y��y�!��A1�T��i���xu��J�V�x+N���x�C���fMY��Y�V"#�T2�ڄ��%�g �Gt�رcY�W]s��}{����#>�r3��� �b��cG��qk�6ۘr���*�F��'nS�{G��a��&�o'��v��d�XjK+EBr�-��:gEݹ�tZ�q�u��V�r��4r_�6�#	(��F�I��E4xᄜ<a���Rkb��!��aؔ�W���>J��in"*,����iѵq��m���T��,N�1kj��bӎ���M�[�v"kl��!�w@�좒#-�
�ۏQ�u�i6c���]�m��@������J���$$�)ʁ%�m�4]V��Z�����aLٖ��Uɕ"�瘉̻��⓵y�@àc��J>@Ġc�H�=\ǉX�YjD�����,�#ts�F�0��/`�bG��D�ZUP�5d�5d$�^�8��d�����(��+v����S��Z.�Z���������j,�����U����*��7m�8�;��)���m��e%[T�mŸB�z��1�ެ`�acL�)��.'��(Rv��v��Ӗ��դҌZ��]��PҶKZݩ��V� ��ED�Ird&J�0+��OP���M*��j[Ȫ�w\|Pt:�)�ݚ&L�h��`�"�dFU��Aǲ-�C���V��7�1��|��A���M���}��o#2AV/p��N㺛�@j�&��-iP=YX�;�6��E�:�H�Q��M��P�j��{J�z0����M���l��ױ{}m�3�g��Y�F{��3�gQ�#>F}��Y���F{��2���g#;�����-4��Vet�U��-Q�D�:�.�"�jڽԵH(�n�\j����7�qm��ȶd5��0ԥV�����w���f�u=�7aw0�o<�v��qA�-S�ףh_��QYٱ<��,X�RR�0�f�Z�v����F�T��eƄ�`�ҙ�Ǌ�V�`Ի���)��-�	c�XO|��:�^vQ�Y���Oi�y7�bJ��9��SmD���M"�l��W��N&i/HЏdy4*�T�����}:���vJƤ��C#Wɐ�e�Sk��/E�ܥ:���R��Y�E�0�Xj�0�?^:M˕��9�NF�xݰ��etY�5ER�rZ���6�.��Y��o#�F$i���=a+��ӾP�ѱg����T���q1����t�$Gë����5Auo]Rkm3XI:Ɍ�)��9���yf��rt@"����v��wp⃣���l�m��kۨm����ѻ}x�kZ\�N�Қ�m��MgbՆ\��;�D^�W'"�	M��uRi��auϥԙ�;�[�{b��I�	etmГ�k7eJ�]��"2D�r��v�р�Z�&�$���
s�!��U��!��pI��4b^ a�F�Y�G+ntre��̏sB�g��b;�BmU�沨[�KT)e��#���|Vq�<���-�r�1NRqc`���*�Սm�u�톅�P��E	[X�3��v{�V��-�:�SF&N=����U�;3Z��Us�gu�r���3�k<Iw�v���98���VQ�ea$�t�/�S��Dv]i��mK�Qn_qD�I�G���Ӑwc��a�M��n�'��|����h��8P��鞾��޺}c�e�g#<��g� ��wm,éT�ߋ\�:�o2UV�]��$���+g,�fk�B������a-|�m:@�XM�='/�`ǭ��EJ�gn�4]�͌M��i:{���7t�H!eȄ�����X{|��.����2
�]rv�[B���a��!ɝ6P�%��HiY_L7}�:N=y��ؠ�m,�w�[5�Ӯ�Kv���oq�0��	p*���C˵���VH-mӇ����eR$��
(�d�ՓkgR���V��hGZ0����Jd»����D���{��}�f����y:<=f���%��b��I����Å�>[և/72�w=B+�ߪa�V�ܷ��<�^5n�J�ț�8�}����u:�4��I��r��������ϯ�IG�aw�B\v���c�M��L�p����JQ�o�s
��lE��os����:@m�P�w�e�O�e�/�-����^<��۷���;�M�_o<$������s�B�����}��a���Uc��y|��G.x5Ts{j��=�_rw�FCB��-�pO[�娍�KC�����:�j�w3�Y|W��˺�}M<{�ʗ
䲻�W/�j���u"��l�Gq��Qy[-t���3���A�4=��7���v��q{�������'��y�yY��f���!�"����E�� �˄�5v�Z�E(��sC��SX���M��9j]��;0ak3v�64�q�Ict �i�2��)d�`�<[ ����2�z�9O��u:Jt I�����R�\�&�zĠxuW;���o#QfW�7�Ua���Yx�6,���%��z����V��=�iG�O�w��]�.����ӸB���}��v�
���زgM��l�qݸU��,�7CŖ�q���Ѻ��� g���Za�GL0�_ $�T ��̅6adC�;[��21n(�����<�q�81�z>�w3ݾJ�F�Sj렐�))$a��ݼޮm�kn�-o3�u�fnffs,���؃�B<y�~�I/$��I,��,�	$�I/n^�u�}�� n���� ��{�t  :   �33����9����Ӯ�t      ��}�    �����<�w��ff��wt;;׾fv�@ x��� �������330�����3��f`737w}f��L��������g`: ����^��}�ރ����  9���  �}��   �33  ﻠ   �n�7m��$�I$�I$�K����d�I$�I$�I$�I{�Ye�I$�I$�7~����ܒI$�I$�I$�I$�I$�I$�I$�~��Iv�rI$�I$�I$�7wsm���l��$�[�Ye�I-�,��$��Yd�Kr�,��I%�{{ym�I�$ fffs30{{{m��e�I$����$�Kr�,�I%�e�Y$�ܲ�m���.�^I! ��vv���y�`C=�u�ff=�wFff`7>�Ϻ���$�I{{{6�,�I%̲�,�InYe�I$�,��$�[���r�InYe�I$�,��$�^�Yd���ݶ�I$�I/$�O�$�I?$�I/RI$�iw$�K����I$��I%�����,�I{�Ye�I/r�,�I%�e�Y$�ܲ�,�Kwv�?{g���d�Kr�,�I%�˗.\�IfYe�I$�,��$�[�Ye����������n�����˖I$�w{�`:}��9Ǽ��^�ܹ}%�]�$��Iy$�~I$�^.��I,�,��$��e�Y$�ܲ�,����ffc�<����^^^I$�I$�I$�\�,��$�2�,�Ir忶�$�^.��I.��I$�I/$�O�$�I9ՖYd�K�ԒI%�]�$��\���$�[�Ye�I-�,��$��Yd�Kr�,�w7��.��ǹ���5˖�l�K�e�Y$�I$�I$�I$�I$�I$�K��m�����33�����Ͷ���˒I$�I$�I$�H6�m�I$�I$�I$�I$�I$�I$�I.[{m�I$�I$�I$�I$�ﾧwRI$�I$�I$�I$�I$�I$�I$�_}�������$�I$�I$�I$�I$�I.��I$�I$�Ie��l�I$�I$�I$�I$�I$�I$�I$�I$�I$��,�����I$�I$�I$�I$�I$�I$�I$�I$�I$�I}}}}l�I$�[�Ye�I$���{�ٻ�s��g�}�3�z�m$����I%T�tǙܶ���;��3=���.�^I ��;����� �}��}�d�I$�A�%�I$�I$�I$�I$�Ym��$�I$�I$�I$�Iho33wwϺw�`A�xvv����}t< {{{}l�,�����:�n�����=<����������}uUR ��"HA<L�8d�nFp�en���
N��}J������4�!���U��T��P��Kj�nv���gte�a�ˌ�Y�Gr��Quu8�^�h�XZ�n�Ц���/r��c�s2n�]T�՚7S\�%�^�T�qUj�U��5��a�{�,�h�LV��/zl���n
�UQ��*lp�sv�c�$���[k��x-[Cx���w)�XZ�_�m�]Q�4�yR���Cl�x��ݻ�I��4��T9i��YI����3{u�gMI|c{�"M��RQex��!}U���:Qp�I�Y��3y`���bv.�O:�AC��X� ��r�u�j�Z�JՏJ�/��Khh�E.���&�c��9�5� v:� e�׉��ҟcvRͨ�%h�<�oYUsv���Ï��B
�ų����u�c�S������Yp;�˙�*��7����N3^j]�.��Y�z�2���}��]g�
؇��ČPu��ԍ^E��
�;��,Rc�(5mJͪ����/F[z�T���ܧi+�q�X�o%u�a����*��O�Q䳊�mt���!�ujՙ��Jz��z��v����&ܛ|'��A�����uW}8�"�j�����U��jb[�yk�_8�Tw:��
Fi��(9vP��Y���{�{�f�@����V��Teռ���V5&�jL���JWJf˪ݴH�/,ݨ��޼�Qt�+��[�+8�7q�T�:�V1Ò���\�3b�$��Uٞ�=���n�x3f��V�lβ0wkRh<]b䖼�Ұ\M��:A@���b�˵F:��	�O^J�x����L�n��i6�\�T+�:��x.�0C5.��`�TQj|�'7�n�>ގ�eI���	�ǭT�:��ʤ�UM�r0Z\�|����Zq��,�l��)]q
�+�݌�{��u�:����s�ed0��[}�����3B�R�[�f���:�ӽN@�i�Q�;���v�Vf��TcMB���jam�H۫tCM`��7�_nEF��[-uS��9�ܔj�p�MNW�;kI�QdX��2�B�r&vTQ6HHӮ|�Ql��蘕�E�/�����Ϻ���k��̹��:�E����0��$[7x�^-�z�����)���ICnAH�9F*�{���F���������L�W�Œ�αEj��L�K��TM��U�V�Ѽ*5���ն֎�,����A�����̭a�R����fؗi.tv��|]fdĜ��1W+V.gvhd��m���i�gڮ��{[G����rWlv�#�J����j[ʅ2���T�*Վ�di9����*�L�H���Z�PD|��B�ή���?�-�x��a�2��ek�/�۫B�Gp�8f]R
�t�.+LBKT�*ѳ5W�V�ja���dU/6��r����Ó>��Q��[r���,ʪ�w"����#�/35�7�pW�&�r�Ŧx�w�^���d`�������o�ζ�'Г���8VmS:FnE���_SZ�{e"��o�d�^V��{p\��9�W^uY�ss--:���/$�-�N!���Q�t�g��!t#nԻ��;�r�Ѩ�2��2YRB
�⼢`��!hk�lu���f��'��gS$�:�xT�I$2@�e�#q7	�e:N�"�q����V���{�����Z�o+���JA�5�Zi��%;|��yrU�[�a���rڥ*�*���ӻ����J�vr*˕9k.|p����W���2���g)gS�.u���̗L�9LVs�s��$N�Wf�0w*�����m�����G4�����)��K��Ry���ł�R
Ҫ�Ib��hY���"�+:�JPF�o,ݦj�ib���T�T���?�-��7j�v7�b����W2�1[j^�6���n��������]����"��R�gfp���T�^�U�Q-y#��N�|*gf���[%�UWQ�l���UK\s��뗸�\N��t�]U�E�P�.d�!7%
�|��^��;P�V����dlwD�ɶ�>�J�!��jM�w�-!�#�e�Ǯ��pJ[R��a�\���ŃeX:�!ɋWº�u�����5��YT���ʊ�#o :���U!��m`�8���{pD8N�)��l+˜^f�H��B������y�ʩ�a��b��v����{�A%���]��G9��}֯Y�Q2@�u5w�f4oF��c���U<Cs��m^�u:�yw|��d���\+.j)��YOcUY�\0m��J��!ǂL��L�ВѱF����e����@۩#�;�Sq��H,��d�P;�֢�s�RS���KV���l׷9kۜ� �Q��ק4Q���[���|*�t��v��j��\f�Kn��151�؂��W49��*;`��S�-`"���e�v�ζ�>9��S�}n�~��7�mٻcKͨx\m��EX�(*J���}U������������2���yoHاy-<ً|쒞��U��ɜ��f��iΒ��6^Ư�5�ܕP��k��c���^��"��U��x�S�9����vvN��^��AM]Qʥ΢ɏ+/;N�;='tA���0��q�]\��2Z��I�ӑ�\;��h���? �:�n�����LȮ���c�˰zhs��pAY4u��5�}�k��:��}�0��y�v9�T�����,%���"���j���;�!噗eWG}ʅ��7cdV�N���u+2��w�@�\��Ʋ��w���9n�u�J�+d�fܜ�_W�nckkIU��Z�����o2F�B��Z��p���Lۗ
c)�9t��V�;ޛ�_�.�Z^@�;	z��*�zH���p���G��Pu�u�v�}n��G\��t�K����h������0kX�W���n%�Ćbn#yū�.0�L�v{NWKk�%���)��f��o��>�T�UVU��H�/��,e[���s�{*��(����b��(L�n��\�H�ǳ�ep�A[׎X�\`�֍��
s������s�3��'SV��������A�M̒��[��w���N,f���C�3d��z��U���uM2�e=�5���ǭ��/aS�As�5m��tm�-Pv��L��.`eWe=q�a��]�b�.%�7�Y��w&O�8��׳�~�'��7b�7WD���D�ƪ��0�:"���oM'���TAu�e��}c�s�iܽ���.)���u9c��.n��y�q}˞D�I6�VJ�z���C�na�\I�����}]ۜ�JǷJ�+�^'����4aRI�R�Ɗ�[����JBu�����[o�+~H�!�)�L�S��I��n�J�,ώ����Z�vE�jވV#!��)�}�tp��*�j��9���u�=S���9f��N�ga��AN���m�@���r|���]c����rݎsBQ��]��.-gY��fH�I#����'B�r��D�K���W^�&?)�ª��� �������u�e=u�dS���p���of��Ax��\��V�����	2��W�����U�|����9o���u��v�'����*6��&d�
��F�Z޶��Sq\,QǔU��G�^��E�vh��ɽ�u�޼0�bو���4�{וM;�+δdk;��+��4��L�3��Y�i�5 ^^T�.2AӵK�:�NJp�c*�w���5�=
�.0֧Af0էU|B�="�]�m�� �α�3�V̒�G_5ڇD�^n��y7
JL��15kyN5�z��{k�`'��	�ݾxA��JB6��G�ʕϊ�A��Φ�I)�:�n��9�c[&����w����b'����m��٩�����)�j>9��wv\��*mtФ��:�m/��T�].�N�j�C`�}�w�WJ}��q�ט[�B�
W��Ȭm��{x��#.�p}{�Q�I�b�y��n�y�͵f`��԰=n8yS��ks9-Ƥ�����c��7!��.��󒃾R��d�4�ֵ0�uwon�r�f�%�.[v;���K\s��	��a�Lӌ�U��οQ%4���+������3*����J��E����9U�ё� ������xk}[�%ǔɺTJ���J�	��(Hu����T�9�z�SƇ(S9.��LX�-(�]m���K׏>�CD)��V�6:��f��Eu�IMXis� �׃�i����
JQ��޶u�ai��Q'qe���T��o�ܥ�
K���`���/���T�}Sm��r&2�";r���;��t3s�{�faC\wX��ݎH;�˹+�+�enTٽM�4��N��	'zG_��;�3�w{��}�,d8�v��].'�d�wh/�fS�m;Q�'1�kTu�O9��K�t��b�K�痵K�yp�#�pP���%��=�h�Q�s/ƕZ���#��_ޠ�v��k��J�P,f�טX�x�9P؏p���L�c���]J�V��@�6��Vn�y[Lr�jY�7E�=7��kg��ή�ʺJ��7���+6�])5r��l��;�˅�*赫Lݫ�	v�$ޫ�.�N�a�zU�Ȕn��w�u�\����{Ƅ|VF��ֽ�(�{�1�}es���c����nv�:'��Ro�u̻��\S�R� ������:&N�oC���/7���6�{��Y�>{2���Y�Ր�<�Jh�\4Q���y�6���V��ӑL�;���3�7�3�k�\��Թ��u�Ĭ2��f=|�i�E���H굪�NTٺ�5d�e���kqn:����Ss�o��tif�};5��������|��ꙹM`�{+f���Ԭ�=�����&��[&���u���5��WBX�ݹR���]�7���J�]3��9�[��K�*��h�{%+�T��]	Z2̧�7��n�Sy]��2N*����.6�0���j��o2t�ow%H�J=-�,�j�T*��G��ˊƍ�2��ّ���mkŮ���%\dg�f�n������|�v�½9�����q�h_k#!>=/q�"����bQum�Q��=���{�t1w)�W�s�һ�۞��k%eI����A.�T�/)�#��.�Í����v�?�����ULQ���zn+vȚQ�g����gV2�3��v`�⋭����F�I�}�1YN� �V��X�X�Ź$��&����Fu�HvU/;�E)xV�f9�t�j�RuB��5fC%��&�;5	r�j]͚ɜ��H�8��)���2��2#��w��X�����\v�y��>uan���<�r���H�U2$�e�!������B�>��u�J9�e���d����L�]*D/j��f�-���ݵ�X�ߖƁ</rqi\�wg�I��\�yZ��e}Nfbr���-kx.�㌖j�����ϝ}���6���ͳl�����<O��;i*L�p�@�=�.�k��ã&����v�.�;옍l�8������C�Y�5��eJ�6�v��W6�e���2榩CN�����f����]�.֊{�m���yǛ�pZ�ԷF���ی;})j��ջt�l6��L��n��Z�^��&2l�Z�Z+q�z���|��Ժ+�oK��y�9��F���&���bU`�����3�=j��)���EM��Y7���=�xw٢d�B�66�˶D��%�Y�r�' �҈�u���,I��i �mzc�.\���EZ��-����&��kF*ņ��R���SQ�d�ư��S'|U�'���::;B�;<ŋ�Ҧ}��r{y�%K��c�yB��3��Ȅ��ηC;v��횰F���_Wl�ܜ��vW2]_C2���2t�aͽ�Se�8�)���z�K��G%L�;o\eI�J1�U���d�������(^�̖5V[*43���}}9��֊!�{.�;�1s��t��oH�(;8{���:�^�;躺�nژu��a�$���[�{��yc�C9
Z���U�	�W;�;8�R��"��m���YD'��݉	]��H۾E��i`�6�dq�Y���c��X��v֋�`��w�#�/)���k��<�-;5�%nN������h��eM���s�*�ަ)^�-o
��R�c���$�$�H�6������N�]m���m���x�u�v������跺쇢�^����/7�7q0M�uRZ���ci���r)n�RԢrl/4GUt9�����C��;S9\�F�%�m�{��Y�K��k�oZaHX�[�`�z�zm���Q��$�C�B-8,��ji5��st4]���u�G�"�ܬ��֡�q�]n\j���P�n퟈�\.S���=;�;l���nՎ��`�-T��Wf�8޵P�ڻ�
�a�W���	�:8�.|�+\������W�Ce΋O$��������U�X�PW�p�o"ha�F������÷+�B��r�r�W/��B3����1�}���Q��1�v�!����P�OUnӱ,>MF'PHDD�a��
Us�nh+n�n"2�gsSs�5��¹Q8�.�T.����fDӏ�S�k^Vّ����E8�8��hJ�q�UҞ_(;�tt��U�/�2�Mgi�zX�{41��{9`5�m����,�mA�����t�
�a�=�IJ�4��(⣮b�y;b��uG�>'%��j3�ʐ��XE���;
����Z�>:ۚ��m��ߦn���H�b�i��莺1�R߬����^ڽ=���̺�z^k��U�G�-J+yh�j���pg#A��3��Rڷ��L�س1�L^�un	i-���Ш�	�����Z&V���5Ë�-���#�k+�Mq"�gD�.�1��V^_�9	�ph�����າ�N!7w+�[9�����E�0�f��Myѕ���Z��U�j5�/&t7c22g\滍��d�+����R��cF�f^���Ù��>����U�y�>�9��3�H�"�z�*Dt��u����ga�vPwG5өb���ƟL�Lq��ޙ�C(��z&�UVÚM#Zclb��KP�����oB��k!���	��Gy�B��*������|˧Ƹ��q�W�Eɍ�T�����D�g���,���Ȣ6>�f��1��Q�I��ï*
oq�5�Ϸ��G��]nJ��A�΋�3{�IUzy��V4+�iH����SŉЇ�,�ă��9�Z��r�y�̛b�Җ]൙H�RY���|�Rh�ʣ�W��eų��:�u&�\"����__[������0��kp�_5����j������=�Tݷy��]��jn��k��l,�.��.WL?:��`�w:���*;�].�����W1:�ؾmÔ������9��{.��ȁu�䬶;4�%�R�*vB5ٸ-	$�˖��8��uϬ�b�[���v�#E��@^�������n1OgP�i�h��l��t�������Eqk�fs}��ͻ�)�\�Z锱c�ڛ{"��Z��K�ݾ���*�f*Ôc��R�X;�et�{Ȣ��E��l�� n@��t�����������ue	M�6�[Ts�y��јs�$m�E�ۜ7y$2�֡��V2�Ǣ4VjY�xM<���W�ƞ�J��|��+h����vP��K=;k9���X`���zAź ��L14�ͷ��Xm��ڷC��+���큋��w>n_f�Յ��LE�v�_�#�;��vpÝ��ʛ��	���=�#-��yʜ�@C��銨[�4]Wip�ŬC����x�3����"fges�5����j�93�V�7��w&,yigLE�4k��tm�Q��@UAE�+�����j�3"�ċାnI6>({��v�3��w9���`�$�����1�v�,�qa��Ъ�n�:{��	:ouc�r��YˍZCx���r��R��q���5Īc�rS{�!�iU�ˊ�t�f���A�f;�۵)��,�Hu�V�}���7��Ln�i]ud�V-������S2V���B����k���w���/_�*u\�E�����27C�7Nn���{�p�R�0���'�����īޕ�beTU��U�
m��%���8�,\����f-E�3B+w�yֱ���N��b�E<��|�Loy.���i�kc��lbڔ��r�]i�C�3&a�Ukc[\V�4��$:46����r��J����jl�^M�s/oUJ��	U5V�E1�Z�T@�g���:��E6	�pv���윙|u��H���}]v�v�Bt��Z��j��6N��c̸���k�Jۉ��#��Ζ-&���ΉzfU[�N�*;}؂��t;�M�N���5BP�k<[cv�z���$����Mմ������}d�����֥<��9>>�Si�==�+����S���L�[�s�xl1Ԕ��F�U�Ą<۪̇Hu�l�Xk�Ju��mU;�'"�
-�N�Et�`%�G�.|��NV�s������5i�Mf�VY���]ۚ�tW����]�Tid�3���'<\�M��{�h(��b�]>��p��Iպ����Gz��v��Y�4(��Rd��_t'�ý{�.'��e���ݓ�͔�V�4N	�vZw��Ĭ���쏦]��m��ss�B�!�xl��kw͙x6���!�(C�ꥤe�-f_��ڏE��,���dn�͑r��o�⦘�Q&d�:UoH¸j$��٦3�K�����@����[X�����D��� ƱD��x���D��n!�8ě�ʢ]�μ���z��X��AiQS�"���T�ce���2���d����ّL[���ksq��p�`���LK�:]��u��hdܾ�}#�d��t&m��V��$���q�#C����{���t��
��*�)Z7m��ԗ�=8N|#�_l��1p�r��u�gcv�]��M�rmcm��}�n�-j��jof]K��4ۼ��8��h�t��[��ii��t���lM
�1���Q��ǻ�[Y��6�+z���0b֔�c����V��O���d2"�l�;�v�Kb�׏��C:��l�X6�x������u��e�Z�+�[i�cM]������{�I%���+]���3�vM	*=���+�Zy+��up4�X,Q,<k3��n���Q��JJ�-�N���k&��|�(6�pj�H9�꺅�6�����ޚy�)���<ePR��\�^��ĥ>��^Jka��=�eX�&I��;�h����9�2v�9Yۼ�x�u�𾍽p�6Ҿ��Ť49��u\�H${Jmf�42N9z���W�;ˊޤ����t�Gv���s����[�Q|4M<�k8�����}�M�y�N5e#L7��^r{w�����]i���J'cUKT��]P�}uɽV۴�6�:���1�UI����{�KT�����]�:�l��J3��P:םiVÙ�Vz�*�?���]��8Lʉ�H��U*�N��y �5���2����&���Q:��ͩ�%�c"7��i*�lB�8��9�h�v�΋5��T
�QJ��Wa��f^i��Y2�3�1!|�p��<�Ph��{��vª�Xh5��M�:��:��2�we&Y�|�uQ�蠊���3i���5G
�3�YWpc���V�Rh"�-����|���4����^��O����*�4�%��9�KZ��׸:�V����f�vwL�v�N�,�=t�`�д�L��$΢��܆�y\�k��)jۚlMe���j�mS��K�,�sZV�c�ޔ����4�܏�U���7)U,J���Z�]���Lܻrd����f�=EGف���cy@As���)pp�4GS��S3H��R��u1^I8d��R�����L��`��v�=u�ڸi���jK�Vul�sk(����ڲ�vl��{J^�.��>�Q�����E��yw���H����{�3�WG��%��Qc��cۋ���"����X`UFӮٔi���0�Ƨm�y�k���8#rl�I�󙙻��퉲��>�!���s��1�7��t��x�����9��;��^j�f��vɩ�FE��}%��ٝF_ˍ<B�8��˷F�\O�j�)�>˵l�U�}��Ua�]u۾�l�*��M�7��#�
3�¢�E�otK�z��Et� 0^�P�����n��7n�շ[*;�Mͪ��wv���E��sis��Z.�\�m[ñ��fl����W���МZ�RP7���쯬���2f>����,�NJ��k0<��u-6;.�iϯ]y³.�P�/;n<���F�UV���	����q�eֳ�lt"u[������[F���δW���{S+)G�+���_*W�f��;w��V>E�o(�Q���zW ��xn��q��ۨyM��J[`�;��|��ݖ�t�2�bTi=��s��*KU��:��X����lm��� ��5��`�U�O�U l�������}n
��4(��P���I�y�u�Lħe��1Z���;t;�'S� �>2��-�L��fY�)҉j8����3
Cej;�N�P;��-*��-�5$�z�!�Yp�Vp���!�}n�\#f�ɺT�;�8�/�	ʏϩ���r�\�y���_4��d��ԭ*����=��x���]ZAf��b�-t�S]N����''�x�qy|����]Z�[�Jh�~�F�wt�s6���.���Z�}�27��;'Ljzj�T��c���]BT��w�u.�9���1���������0�����Y�0͈�����3f|���[f;��Y�}�9����"	7���/<�� ��:���iͶ��o}�,��I-�}}m����[$�@�A�wI�ѣ�� �"Fa�ݛ�$�@��Â0`�$����m�Ie�m�I?}��:����$�^��I$�I/m���z�3�����^�����3� �Ԓ���N;��.������!�`�s89�uS�nf����ʪ�U��\⸩'F,%���6H&�`��1�%�ڼ���%���P�b�	5�&k����縶�w�p^�e��鷔v�7�2��T�$�]^��;"����䅼�Ǭ�Zل����8��!�]u׎��|��􋸶��j�g)�l7|湏�T�����rFJr��p_lWgc
���9�.���vڜ�nt:�x���w"bq;�jf�S�Ms��6Ĉ�D� ��3�$��Sv��5���g�jcmgT��]{���ro�������T+�6Ћ�P�j��qToS)��Yǚڳ�U�����5o-��we��RU�N���F�M*�wY��.�]c]$�o�;������w���!5�T�YQr��^Bn�̿v�-V�쵞�eo���*}_w��-��9I�T��6�~Tw��R'��4i�sB:�,��QX�ʩ�b�l�j�.���u��H�Hop�\=��kqv�ח�Ц;�,�hU#]�=�ڧ-'��&4s��Vr��X��.�2�S�  bc�	.rڳF�y��	՛�ݢ�*};[7��3܇���ǧ���v�f�V��J&�IO���wv�LB,��@�D�:ĞGn�;u��'I+(I΅�C��H�YQ��y,+v��vQ�PNy�W�Ɠ�9/3"�7UA_��^^���F'{��t�DJ��^�	��0��-ī%HҬ4�۩EI�g>r��Sy�Խn1�Ɍ�&5Cl%{Jr�}�Ħa�c]u�L x�PKЃm�KjRY8�횭[-��z� ��?a<�{�}�+������V}���uyV����f�b�Z���&HWƎj�A)�Q��u��3�Fʏ��d/�[�2��Y��~۬�ޡC$�dmv�Ec�n�E��=����K3� �RGWZ��R+{����WmL����.�}VK�d����bZ�T(��)5B��V���V��U�.�
X���7�K�Fl�i7-[�s�ġhTpe�"��e�-qw�P�^��!�Q
QV��8�=]k��n�6��L"�ї-�e�u���a�J���W`��4�r$Y�I�B�Y��^���P�ǀ�btqr�
x2m"�Ý�%n� �O�t�A�;��:q<ڸ�[��Џ����M��uÐ��մ�ږ���c���[.��]�5к;��g���4�>� I�Q����(�v�i���)���ü�:��G,:���'ɺ�'�;��X|�L!�Ö���n��P���,��0�>���?��������陔`�&'(��j���!��A���D=��`��0�KB �D"��e9�&����$v(L�iBE��ءC��{�^���mzA���,qǑD�v���B5���g�X�˜g�l��F��s�Љ��m����B>,�5iʣ��4@X�+�#�P���]CB���<9}T#E���K�rl�ٸ���<`;P�Y�xq�,��G4�G���,�P���smD�P�{���ߗ7���lCr��� /�R�G~^�����4��e����s�b������*Ռ��A����c:[��q=�E��:���y��]�+5���cI#\�uΛw�h��W���Ո��}�8���6Fw[y|�ո�����o������n����\=�J�s��^C��u*�O�P�&J�X9$�a��"�h�>�/��v�z��BdAEG�-$��|���в���|��OŎ;zS� �O�i(@�g�$��};^ ����B�aP 0}��"`PP�Y�N[}�x�4�����HoYpJi4k0���vJ����$�(E�$B ��	��ǇcX.+��zS4S7� �(H�NL9�C�#Y���L��^��� q���D�v�
��A��,����ݯ�&r�$����AI�,z"c�!I�5�~ �<ˤ��9��Y"&�!�
��C{���#����:�"���$B�G�>�9L?jf���)Ҷ(�~�	�Hr�z���mt�W~ǯҽDh�Ѥ1��
�'zӛt�r��;��1G�:�<���d�w��]K����&�&�P{Z�S���3��U_[�Ť�tΏ&-D��Q�RgUwn^B���垹��o}9�9��'��Ull�U�`�`�G������(�F�_�Uf}�UU5�x&�C���<8�.$�� �k5��͚����D�'�yh�����b�'|�&>0��(rHEX�i¡&q2,�½$���R�˸"
A�� 1dy�a� �����՛�h�uQⲄY�4� p��}�0�4�+O:�{j��Ђ�l�G���NQ��FVD�eM|�@;X�;n��>��k����تf���D���8L�&�0LH�f�l���n����M������s�P�\@��1{՜�%�z��W��W����j�{�8���w<�x*\e-h��{��1�L�Ce�>|��8+Hmdf�h��a�4 ��4X��$l��-{w�����w��m�}I�t�Hv��ɝ���n���y�u���C�ޅ�>`���H �h��@D�
 Y�(��3G�@�`I��#�zW�`�.
�� �d{�ޖ��OI%��4"E0��A`�8��|�.�ə#~�,�DM�F��|;]�%0�=&���)/����� 7\���(!���Gu��l0~����`;���� �X��G������e)!��T�YA�X��xrH�mVG�#���(1�4�|��4��5�>���4�kG�`9!�v,2?n|�{��'����S�!��4�8Y��z1ʪ D�Օ�y�ع��o�1H�\��ʤ�41~"��4�Z�}h|>�UAb�>#�[�b�?��4=(1���v��L�����T!K�8ok2��{D�ɭH��m>}c�xhcFU

���!�v�%�������uW&�1���of�ݬ�̾�X��189LZ���D �'u'�몒%R�6HF�-LBR���d4��+��^$IÅ�$",�����U'�,h^��ya�,E�Y�x�d����fH�v�&S�c�&$L�|}'��Yc��+��o��`�(`�Ф�!�"գ|af�L���Zr�(=4">>�K��<���5��e��Yi��P-z#ęX���J'Y���{�C���\~��1hXB
M"A&��5�7��&�����#iWEA:=(N#��A[�.�U1�H��G�$���=��$>
E�]�%G٨��]��j��>( ɱH���L*����v��ޥIު��9f���P�Ć A�?iH!�ꥪK�u:3K���)���Ztўx5jߝׯa���<~~=�b�n8��Jͯ_y.t��B��ѡ��b\�6�ԏjV8e����mU�uS����A��A��h�b��&�q��6Y����%![�����͗TA !"�|ߛ���y����j�r�|R �v�H�
H+� À�}�G
����E�u�������1ho[YTB z@�6p�}��eT�������=iʄ��ш��e˸��}K�9�M��ȄFP�f0ܻĖ������ǡ��4�<=O��B~c'�����B�+�@��p9��{�E7S-�G� Di�|\/�x)!�*�F�����1�MEmb�OT|Y(� ��A���Q���/�5�p��ib�*�d{@˗<f�a�%�T=(T��P�ኳ����uc+�_�<ޠ>�!������r����@�kى��L����=��ʼ�j�p�����
��A�S9K�f[��,�0�ڏ=ט�wfb�ǜ�WqU��I�<0���|�˛P�R�sC�>�䈈p,�$�C5	��$4�Z�1@Ah�h(��
�V
d�P�����c�����H��cW�@�a�!Q��_� ����~qT��!nq�JAB���w���r*T䏤R�xP&�O�i�6�}M���d^�;�)`D]���[ǤB2u��ȃ=��W7Y<R{,��eBv��z�4b+���ک�'�c�!�%�@��C�����,|,H�G��c�&�E��Îx�hù�|G��@�"��0X��V6�0���]K��	��U�$W��~�e����v�i%���I�����#��+��7ya�w��G�i^a��l.���9�1A,xOA<�Å
73n��/�La+�e��JU.M�ý�f8��G��O����fsp�ͦ,p3�fD|XE6��j������J��d�� Y�P�^@���/u�҂FeA��j��z�Œ��#�	<>�������Q�� �&0@����|>x0�?w�4�p(o
�@�!�'Ï%�K�Ó���QZH�C�O�L�x`"B{U1%�9�a���YL��8��!3�������!�&3�������LW�P��&�!+KH ��l���,P{@����w�Q�-�@��A��M�w_�{[U��0���Bv���-�і�L���<U�]��<Ac  ���*h_S4W�levd��,�Wd��|�_�䱇����U;�q �H��"���|HI��Cro��V�5�P��8@�N��@��+tw�u���|��u�uZuG;sg�2�Z�rY�HJ�Z�64dQ�j����̛D�ts*
֘/��=	/�$#��H.�|�h6�A�T��E[�~�z�oP>0d='%�s�}Cд
��Qn���-�D8�X�S�|P\Ј �Y���,�u�g�q�$B��!�R&�"�>�f̬�g6,�������D�i�Yo�x���C�Q���K�;�����V0p�< ��G�y��n͡�@�(Rm��0����Oo��u?fL͋%!B�b��( ٱr�"IP9���z
Il#EB�3�i���ם��߾�����)�AȤ�'0|B�0{�V�}訩�*� �|�@h��	|:�����OY�����E�u-	��Ob$�UGz��Eb�>�q�ّ��������^���(P^1!��*ߨÓ��@�^��ItXz����s��:�tP��V�-�^���T��s5�q�q� �A��5K���Nm�*8�-�81_h�#qAIC�~�,���qT��p�� ���\qϏM�X�4�f���{�>0No|��4S��2�Q�QLxr0���J�>��PzDC�@��b��&7<*^��P\Ј ���.���߲�]��9���C�8
�A&gtׇ��9�#�ogŔ���0�M��P#�ǧFhϷ�D�����)5QPI��"�N#I�ȸ��V�b�,B���Is�E����n�C�|�Z��A��,������cG B�>��/� S�ؒ�3j���W�@u3~��N�0E;�r�Ar�YF�j{~�ނ9X�����N���m�yG�f��շ�r*��s��[v�;V�Jn��Ҫ��/qo�W�����w7�n��C�*��}��z�%��^Ą���&{�	Ʃ�9"p"���	� �	�Q-���`җ�'O[u�W��y�����y���f?;W�m؆p�u�����_J�UZ[�t{KY�U�:E�]N����wԌ\�y�n�k���u.��5�z�x�Ak���^�����Ȅ�^�__����'�V�u�W8O����~t-�����Z��!U��)���yW2��ne+��hk��p	�E�ۡ�%fF>�%�Փ۞\��b�.S�e���>�J���D�ѫۗӟ�7*��=���{V�|�+uW#��S�/e'����)_L��j����N��ײ��|� �ޅ��n�0�}��Ovw�{��!�77×y�l�Om�!Z�.v�[�U�\��~��{��,��Ʊ�wcs'&��M�9��D9�@��.f.��&+Ը��5����ie�T�DVi+*�*�݂�����Җ�c��f��P�^t�գn���M�}G��Ny�אZ*��D�I�4z@��ww@: �������>���.\�I%�ܹr��}r�ͷsy�37wW����I$�Ir��$��m��$�_m�ۗ}s�uw//$�iw$�K��I$�I,��r��/m��%�ԒI$�9um��$�Km��d�I$����<�]�K;���Is}��[�����˭InzH�>�v��wwl��q���Uu��}�_M�ۮefv�i&*�IR�Ϲ�����{z�g"/7�㓾s�������w��o�/��8D��w*���DTy��m�<�wG�0���׎(�.÷%�؁`�k�}���<M*E�����/x͍nU,W�^��.�ŮӸ����;dO�{'H9Ӓ7F!�K�f���G<wZ��ٲ�Je��pr�|��֍Ӛ�rƍ�;����:� ���ӓ�Бn��\s`]����c�W��x�ެeft�Yқ����r��!��
���M5:��������fG.���+��j$��tLꃳx�ȕP���8�\y]��)��nVžtJ]��n��%:nN�/��,�cn��n�ޚ��E���#�,�ʎ�څ��YP�W����۝��d��*�]v�$wqj)"\�����)�}�tf����S���vnI�]<܎�P}�d����6����rL�[7����Cv(zL6����ζIN	סFb��X��9j�ed�f�.���F�r�n:E3����Av�X�{(awfؠJ��u����=ZE�"���l⪱Y�KP&�LΨɧ"D*Fb����5{SE��+�PꐌV:�<���
��l.�F��1;�'q[ۼ�r<XFP��L��	Ŧ��֩t�tY:/�Ѯ��{-aJ�������*dbʂܣ����&>��Z�-�|��\ZIX���Gn��P��u�.��X��\��DE����+y�Ri�
�Y�A�c�D��s�$�a�劎gbr�VQ�cE��۰M����E�9��c�jp캻�(��X.Ŭ�8�!,�O&��,�Q�V��p>x�f嵖XW7٤��Bѻ��i�=���	��s�m��[�P���KU֖:3ZT(�ٗG4�ޔ���-*��4M�R3���w��,]�Z2��/lH6
�W�#s�@�Ydur=}T-�ѥ�6����U͵��.y�ͽHWlٹ�0�<3�Q��U��y���I��mq�\Lfu
	��v�h:<tyՒ�L��3���5��4�Tn�Nm���p�@� �A�XE��id�]���Q]72nK�Ƭ����k�j����&*�Z�@k����=���Q�^$��DP6q0�I��[.�)A�����E�dҧ�Z&fJ�cɂ�7'��6�?�{[r<M�g�g&�t�,���v���7�9c�f����?u��f���K��M[=-���]q�8���:a�@:`�݆B2��ݽz����ߟg�{M�=�}���)�"G�������V����gv;5�&	4!��K�}������|�$v��Ӎ�~N�ն�˛u����뇻I�X��3_�U�D��`$�|&B���c��n���1��n���:[���O�q�a�x�9m�~��ⳫЖ�fe>�8��rS| bXw����>8�����Θd B0M�m�H!Z�����ފ�Ȉ��&a��38�|K�LX���-�c��۞�q�:����l�~0}�DG<����hp���*L�Y�e=,���~�����ro��n���g?3wݟkj^`��H:巵��I�8����sl�1;��X�	��qRF��w�wg����"�t�$4��DP��� ��3���շ|p��?���w��I �3���=�-Aiy�.s�B�a�E[Ÿ���kC��BȼTG����_`䑘��9!�e�,X�1���'b

(v�6\5��h\�y�w������:�"�[ݛ�6f_YޥY�0��9La�寕e�A��4?�y3i QI��T�m�CT�t��E��#۹+����@��CKj�sz��iώ<Z[u<M�a�xM�@�n>�'�TS��8����g^�GſS�X�c	��8�&4����������v�����I���KzOws{F��l��~'�w�Vym՟0�#��Z��t����������c���s���]�~^Lژ�v�R8�q739���D�x�<;��q3$5���4~ p�۫oŷ,��&���߉�Ԙ9��,�����&���fP��oo\�����_9�Sw�,D��&V!�D�	��/�>߻6����Xd#�7�3��E�E��6�C�.Sl�>-��rFܞ ΀�32�h����ݎ<������o��m��۾a�N��6ω�w��Ŷ��oI��3&r\�5�!7���>*&����1����X<N|q�Ζv���d��|[�n���Okm�����{{K�fffp3�q3K������z_;s�q�n�����*��4M�kz�����ԣn� ��j&]�U����<WŽx���%����c�h_��y:�_�]�/í�y,`c�D �F2���cEG�9��v�fZ�37z�j���-JM������̝wQs�re)}V�����ZW��[�W�5�A"H�% n�䓫���e3��h}WLu����8}��D{S�Ǥ���~=���ɿ8:�Kvg8xM	�:�oG�~�	LJ��rm'�G�<�[�����:���>���8��x��mF�oaǳwc#n��,0�0DP����n�����7V���'>'����,�Z�V�t����޸���=}|Y�E��ft3i�JfI��?Þ-:�V�l�:M�����8�T��îf>�ǯ�"e٠��S4�6�&�3B0L�"R��4"���ue�1�d�G��x�Q=�V��#�I�<���n[���I�|���|u7�ugŷ'n����Ӛ&���N��������k8"fti]8�������ͫ'�m�볱BLA.jfq�ˬ�=�AT/{r7���������x�垜���G��O.��<GVj�������LL�}�F	���<�i@x�������./S��&�q���V̄xM�;!�|�1����+^�fe�;��@W��!X���%�Ic�����,I�u?��ͽL�1��_�/ٝo�_%��h>�kw){W�u^��ex|a7�"8Ԅ�+5���?C�vOlc���=Y���� a�7�
���[8�	������/"ޥ����25�K��\�����UPq�����	��C3-Q�e�m�����g�c�8`C/��i/y�<π�}�N��7��wќ�M��ޓ�naŸ���x�۩&}�0�Bዃ����|�'D��Le�96H��~��nl��^CQ�1Ν����׮?,�}�_o��{������a�1 txO������nGi�/ɷ.���K0ZX;1��&g\�^^�鬷��<̜v����c�g_8B��r#D�;:���{�#�L[��q9GW�7C�'�U�0�SR���N'J{s�[���R��c�����8���d�;�a>��9��;a������*��(΄����(rȁBF��B���	��Q3zQ��Ԓ�>s����G�BP=PH�*Ÿ)
~��AD��:�S��uC�|QvK�j�z*&>'�{�X�u�\q�x�]�jbf�3�!I��Hf;2H�h�(q�	�8��L�4�+�:gW	��s��p������?a>��_m�Og��PX~~��hD�՚��(��|Vz�w�����,P��"�I[q<�֑ܻ��ز�E���ۮu���ŕӶuauԹ��:�����=2���:7l����"JL��52G��b&5ߜ{�b���xq�xLΤwl��~><�zǉ�V�GHd�i;e��`��G�<D�3Z[�4/`�7�&Ia��D�&p����>��o��-c�]������ ��Ba���}H@�8�:�0#��;c�"fl1؅E;<ģ���oIU���đ"f|�tI�C3�O�b0ʩ@!���K��&�����Z�ft4|.�f�.��C3�P�8�|OE���a���л�����FL�8ï��8`�|X;3e=����q�O͆�N�����.�ڰ�03:�]��In38�u��r�m�;Y�����Ë�6���7^(ߏ��ta��N3>�{~����wx��[�6���%�q�rݙ������A蚯��|sl�s����_[5lS���O���/;1e�� (�,���y�{UMoX�s��ІD�����Zg��hv�@��vpAL�ۿY���8�y>Xh���l\S!�<�iW���'�i��GHD 7;����eU8�d�UC{Q���bA ��NݓF�(	5ƍ�:@�+6���y�n*iN����*I�n �k�%��2��J��V��|��͡UW�֔j��ƚ�Cq��(��æ��tG�z�b{. ���$����O�a�������a,�DjhX=,������X�@�B�Nf��J�}�V]��M�q�G;��C�����N��0�D�8�Ru�M��z��
�h$�gT;�!"���H� ��Ma4���J���Qe���}c�$�X�"����qͫ��M
�8Bb�NW|{���0��i�3��è��8��q�L��h x4�N�
����b����tQ�D���uT��
��d�	����a�鸪3{��ǺK��q��b!X���mÓ?0�ɓ�&�(��rgS��>Ń�Oc���8��cۮ;�=�f���}�Zc~��^��;�$D9���cT,�lߣ�l�sՓ�مTUy�"�o��\@�dx���mJ�"�_ܫ�LI����R�S|�� ���"6�[���8Ҧ���M�6^wiW��P(ګ�ɍ��ݕ��.��KJް��'h/����i�����5y�a�*�&�]�Z�t�3�}6&d���O�aE"�	q)$�|S؋�!��C���\�E%�wq�|�.q�'�۞˘�OG��.X�Rq��^Ǻ� �Α��f���Z|h� ���`�u'3c�L����^e�)�Na��UL���;��I��.TG���L���,����Y<C��N�M�����wK�����u]��-e�16�$��DT���	��*���բ����a��G��:MF'lܕ��«,D�.s$_׸��s/.���dH�C��UѤ=ڈ,���!=�q�g8��S>fc�8�'q<�xȢ�������'C��+����%�T!�J�EWĸ*�`�&
����}u��Y5q���|J�.@~<]�LiGù"jC��,yeU?��*gzl]Մ'Xe�VAU<px���gy�<a�Ѹ0Tm�N��ía�OW^3L�}����r�9�)\�]��.����5]4��n�;t���nE-	!���ˡUO$jU�|Qz��(U���Lv�|���P��ʲ�rOP�r^����>0�	��`��,���{ґx�p�>xRR\>�-5���8�?�Ȅi�YC�(���0�Us6i�}�:m��������F��;�����z�.,�~?;����\�z��h���c�#�c�#�j\@2��-�bT�vfj8�$����fqx�0�'\��ha���g#Ɂ�p&�fiDn>'��$��D|C��h\����.7�F�U�`p��l-��O�0C��$��$r�-1�0�����iꪼ�0��Cq?�0��΀M�<i�V�$�v� 
�y�����<&>98�#ø�a�q=;�w��B4���so���~����4t�pi�=����+
��B�������=�v��YJ\<x����*�St`�-�8|���2;k�}_-�ω>��c��zYA�"�0M����LՍ���S��{��Ds_6�☏w�VdT
�ȳ�Z�0��a�ٴ�U�%��%�ۧL��L߬�X�ɲ���7�Z$�����FUJ�x��A]|�-�>(�a������3���:���*=U}U���:�"~�!�>;�ϒ]3o~f�z�*�pT;�_u=�X?4��D��+c����i��~�!�w�(D�/B}w�PF�Y��Bߣ�}V��3���H�a]�����JB#Iz�3O6�B=���� x���L=��݄�����Έ$�O^��y�v	0y9�#cypw>4ڲݒD4��e>�|E}�o�Ρ��lXlD,$�@�?X �[��\��q�,cO�$�OՄ>�JM%�ǅe� U�to�nW^f9�Au_�$ Ѷ�VօB�'�C�����6q��|�����N�g��\[�pi��w��鱼�i
�����7����Wط#4cG�a�,p� �Ac�ot��v�ڦ��v��w�]��۵�r�CL�:���kə���Lͭ��/-f��#��Ɯj��ջA(���p"19�7�m��h�E}gى#�%A;N˙���G�EJ���}hD�'��Gg����*�t�+7#���N1�0���+O�*�0K�<��ZmG���o�ntw��nph�!��A�')d:���'l�1'��.�~f���� ��Vd:$�D�VC��QF�n�0��˰@���xw@�Ï�Wi`�L�9�z�b ���"������FЉr^���T��~,2��~����Z��s'X�I$�Ey/����F��'��?0e��䙅+$4����Q�gTՐ�;��8��1�����w�k������vI�Nס��֌�~���Z�x�9�柳��Fr��t�.�\P�%[涸c����	v�ʊvJ���qi���bV��c�TS��^�i�]V��ml��;m��v��8[��W����x��'�~7ג�+�94��+Ai��U��Bj�h�0�.8b{��{������ӏ��)�dyV޶:�ҽ�k�{�Xe����XM���;m�;�:[T)��">�z��Y��7׵�빓�^��32e�������t5zw�h~�s�=��}����u�V�
/ە�����[�׳���u�Jެ���:��n2uwN�����7��M�-~����R��u�A�t}XY!���+��|D�L[AͮRq��@��'�o9]���#UI�^i���w���S�}�3�������ۥ��u3�7]b����_!Q�{���s�,u�Y�A}�ե�?V�Xc!b��3x���.;�޳�3c�X͔o]�/���$�Q/|���o��x%Ug]����xZ�����{�5O~<�r�K�]�_�������.�S��-j�����ڃ��1��(�꧊�n��п�Yʥ�}'���VW���#��yx�qԲ�p��E���"�ٗg��zD{ݚ[�I�q�Ò�U
%|��.��7�ןĀ����9��]�C�@g>�G6�o-���\�r�I$�}m��/�����I.����I/���v]�����^�Yd�����s}������m�I$���{m�I%�-��$����uuwe�I$�I,�I$�^�}m��0uԍ��_____J!t��b�n㝙�pu�s�ْ�r���Y���\�aʩ�z���ϴ�T�I�f��':Qu��t�h�zn�i�B����؅�Q챵�E+��
϶�	�Jwg(.$�Mq���*-}f���M[�飄�O7[7�d=i����=��W���jq�q���%}B�i�"�������R�`���t�}��\Z��,�f\�Q��]^b@ңI�t���q���(J�aq�����|:��I�QunS�dn�}�����L��$��X��lSX�[�#�g�7b�aΑ����[��٣V���t\\���I�n�z99�IZ�%ZE
U�X��|ٴ��QBґ��}�f$N>������j��J�����q��9��k^ܖ�!������.�jF�5� �Ǆ��F�mu�䄚����d�0X��'�h|nM��4�&s��]��e�9���l�M|.5�Mց���ĵ}-������RW;�q|�є�jҕ���]�7�w��;K���hBs� �U;k��F�)�-�vxإvZ�Э�5���=�]>F��V�=�Ѥ<�n��Uwz�ێ�f���fY�ê�t����,�w�*Ż���FT�Hv�}� �j!�Q�J}
���g0�ϔ�w��O�
Av�GT�~o�k�\���f�N��ac	��*�Q�tkE�u�*�f�v��_b�ZL��D!&7nV�M��ifw5uip��������seU-�:N���Յ�h�[����u�y�Q�͌뺮A�쁌���&����S1��9�WUngM�w��ؽJUN��X��ڧ�h��j�,���XځҰ��Z���le�u2
�Tf��o ��5�k%�m���1�R�!T�B�W56���/��[J�^��E ����z�A�d�i�����2������7�L�XjޮyO*N�Z*[Ц�Aτ��A�n�Y{R��;�ϗ���nLv��fP��T�W:��v�a�ݽ�)�ٟS��4�|��W�����6�%�@��pyi�M�D���wR�֢�J.pu䩘 ;�[�t�Bű%<�N�i�s�)
�s,*ٵ�|h� �l�m��R�P���%��QoO����/w���PpK�G�����	�X Ե���p�_g��"���d>��JM%���YqEQ��&��q��ߪf}�{GrO��p���q>%�Oc�}F�g���;���ox�<nZH�4IC�O�x����d�~����,�9aX��HË�M��4'�np�w.�����φ���
�ඁm]-@�3�v銺���4|�J0�z��C����B�"��ȃ���>��=Ov���и4D@�'U�����8~�sͿ_�<F,Ac�a�+��x&Y�8�Qd9c��|�Tc�{��G��$|'>w*�x�ʒ�rGv��"��5
��o�[~�|?ve���c�j�ʏ�a3%��gH$Yؼ0�@�h���;����Z���7�E��K}����1<b�6jI:���yN��tK茭][�����t��e�HS�G�b��23��[��jȊʇ����|��V�#H�W�˦XGA;��^��ʆ
��t B�*�P(4h����O�hԧܴ�(��0�
�,�$w$~<I"���ɳ}S�5�P#Ĝ]qC�hh��K�H$�+>�=�:,�ϱ�0z r�0��K} �&'h��o����]O�2d�x��IX�+.
*��$��L�@��a��$�dq?�������đbr�q4�q�2;/�x�����⣂AP��Ax�-�*(|1�#�ﳺv���e�;I.�%��A���7	G��0a�n������cC��G��� ����!vd5�i9Gu�x�U=F�: �$�(�x�(��R`�Ǣ�.1?^/��T<��������q_ ΐ'�_cP���B�5m*L��yP�9��>ܙ����J)��
.��̷��veA�5]z�[�x��q7�������%�O�ax��kx��]v��+��WrĽ&zX`�|O�T[!��S�5h�EPM�R�;wy2�D�Q��h ���䍄N$�E�4x�/�ꢀ��W�t!<,�O���ܑ��"H�9���(Ga��n��	0�ʒ�rGv�㉲��5�0�n��f�f`�-8��E	��`��g��f(��N+��܃~��E�L���ܑ�8�,E��9.sƛ\g�҉�y��섛��r��rˈ%��@�F+�q_}�q�U]!f�@���!T�� �&<Nф9��'	�x����u�EE�����e�EQ��I�&��'���s��}L��Z���A�|I',w@9��Y�bG3dh��N�����4� ���;�x�����;�;|A���s�҉����NX�ϔ�{��xs^�x�?�|�=r�}��@8&��}Smj�k���f��p���(`����4t�E]�3]!�۷*����lu����P�"O�A�k��ׯf��I.�̢&�l	0i-5#*�:, h�A!6A��Z��A��>ڏ:�����{�̄qd8�@x��Y�J>>�*�0H�K�}���K��x��C�B�t?×ja���r�=�s1~�V}(l>#���QT9z����I�xx�����ٙTт���8��AG�x��;�0sOb�8�>�sz*'" ���g��Qd9c�h�$>�Gr�o򁳦���ŐeIc�#�Iǉ��.|;�R�}��ml;�>�؜��E�)��=�#1D4�g�*hъ/7}���>����v�qC�%d�b.!�pC�xڲ�dp��{�b�"q��(������	uG�A#���������_�v\�xBž�M�'�a`�I)4|H�c���a{7#�;6���X���Ci	������S�df��
8k�0�T(�{$�Y�,xZ�<m8`c��ʻ�F`a��D���[iX}���]�4�5*Y7e�I3ҳ0��܂-���'Zk�K��"f:�S!����IF/Aq�DB,�� �n�p��04�bnʌ&ǃ>B�Ls��t��'��!�b�B�����B��x�7�˛I��g?	���a���iȑ�r	�h8�|蘉��8�B$zNh�H��&�5��0�����&�Z$a9fa(��AVX��G,rHs�l�9�߻6��UI��|!R?U)�����{ t@|F�?0���AI<3F/�*cDb���>�:�"~���f�_z=J�iz��1x�⬑�;8���l����������������g�j�!��>!PI'>w*�iF�s�����0w0wm>8�`��s�r�$z��z�׳*�s��G+&��v�JÃ(+@����ǹ�g���{(��x#����'Z8}Eb<��,�Auz.��ջ�_z�7�/����	���H�Q���}V�q��Go�D�2�vUf:�c���깚��c�A���F�A<���RE����%�}�x�[���$e<�3O�wd}uU� �z!�pC�&���k@a;G3������.�ěƟD��� ��X�@�Üz�T����<�/�0�q��C�;�JMH���V\��^�u�%L�C5��i$�ù#�a��OEßEH�'I��߷�z�3>�}��.$w@9�Yt$"ӑ#���;#�����04��#����;�;i�d�C�7�/O_ނc*�����{	G��
��L9c�C���ЄLw�wն�𼼵j�3�0�a�r�=�: >#Ilx-�ai��TC�Ad�C��èB'h�q5R��)\_<�t�(>C����0�.�#�e�s��-���}�&����>�����g��z��v>����!�O�A�|E.7e�R��h���@ �X` ��cn^ ��F�����ɼɝ��ztk��uś8�μQ<�n7|r��p�f����ǁ&4�g"l�H$�U���G�$u�66ͷGSt+��E%�HD<S����#I)�i�{M��n��`�8Y@`�=V		($ �(w9���߽5��^^k8�{�Y��ù%!��Br�q9��fפx��_�f��]���8��Mc�C�qH�#�����uy�324�Z�x�`��ě	��1�Gl�����?�wRfqn�� ��X�@�i�R[�Q0�xᵾ4��K��_�!��%&���x�QO�I$�5���ߝb��4^(wo�.�S�p����br�s�k���=�ت��YQ�.��Zr$|�}C�$w �8c�$���椏	�������K!Ă'ۆ�K��Ȉ�H,������G,rHq9����;꾉�[i��PL�ÂG��{�<���'�g~>�0�u8�����ӧ��RV ���f����a
d�x�f,xxR!�1B0��颵.�u|n�T>U\�����ڏ��r]��C���Q��n�*������?uri�1�A!���q�KĒ�a�@^���^�Sz���+u)�{�˪h�*�,@Βm�+�s��k��h�}B� ��<H�c�o�T�A0�|zo���U}w|�.$| t�cPO�\8��AD�/8���s�2�-~�F�a�Yt!<�,��YX�s?�{�]oD�fc8���i���T��
> �(w wl<q<��ĕ��=�싫p��>�4w$�",��NP�#ÊC	�l�j�ea�̺l=j!�F9SC���ďb.!�`�/�������qDɃ��74�=�K�4�$~=�����U_]=��x8�4�T[�Q0�i��C�1����5v�Y��9����G�e�S��I&K�Y����)Qg���)��s�ܢ���C؜��M��[o���Y�'潡���e����L���r��
� �5#S�5�;�Wڬ�,z�=�x`���J-�¤�kJ�D��\.P��\M������ob5���L����MM�剸���#k�;t�@h-,�k�wp�5�U�x�+*�E��6|I&�����x˛�%�e�]B5;D�!���#�jD�I�c	����R6�UM4�J���&�,�O�V�|C�W�,���D9c�C�FB2S�R�m<q9G3�_c�d�UZc³��ď�<�QRA&J��%���ޭ�e����:j1�	�&�PQ&�GC������_z�e��$�.�#�e�s�}E���B��9��ܩ:"j#Y�D�A$�L�;�;�x�8�%�`��gY�����i�JH�'(w�iF��Q�Y�o��^[�]�i;�A`B����E���ag�I���m&��h�Ě�I�:�. �T|D8�wo�9�E�2�rJ@w��܉����Z��>��X>>��i�'ò�7�2l_�`�4A@����4ĪP�*�%d���6��ӵ[�\�W*�\
��h��lp�:w���i�����
Ŝ�;`�l�B��B������$"��"2�3ڍڽ�� P�8��3�*�| z��Vф9��'0cӚx������K��g������)��I&K��ƛb)��cj�#�30̕�;�|�O=����8�8�.Ďu{�/��wg��y�Ä9;Ax�pc�!H`h@����]~��V����?�Y�ǈq ���~�N9�M"`��>�ɋ蹪��9D8�It!%>�U)����=�p����UL�������z<� ���>&J�7s6Yޕ�/;>��X?�9I�T��KĎ"�q0��vs7�~��ꦩ�������Q9E����$�5�Hяq����9�A2P�@��x�l��T�a[�rN�����]���+ �޷R�����
�9���K=>䷂a������:c���c�s�����#tۼ�2�Ia���JȲ�s���\�y\���a]����h[����,dE5�s{�\/:z�����܇�oQ�U��N/9�������7������v��ofi�k��q׹�.�;m�*���˭��嚑�&�e���[u�ڮ�P�1x#�>e��c�{�PuEý����=r�@jw�f5�v�WC�����s�����8���'n>5z^7vTW�yh�ԷKW�<~�	�v��ͧ��G8Ѯ�XvY:.�KV��9�o'��n�\��\ާq��ߩ�ǹ��,͎��K�Ό�f��}=��zˤ}��vz�w�ߥf�_�}�RZ���;T��#�|�����w��J�y�B�޼UJM�6%�S;���/��~����΂��Y��x��3��X�<���Yf�R^�B��˜��/��IEVL�Y8+�禼ꜱ�m���^	�>u��I�|��2̨��^���ykz�}�鞱~/�b���ޮE�n;���^�6���i�pCI�r������2�ο<K�w�iu�
��gc���$,������?�={��u��%'�h/}�^��{�7�<Ͼ��  ���7www@��\�r�@�x0I7R�Ñ+�,Ĥ��a�I$���m�I%��m�I%��\���]���$�I??9fe�I$�Iswu˖�l��m��,���,�I%�-��$�Im��l�I$��fg~gw�����[�s����T�%̂�w��3�m`~�ڧ���ś�2�n��J>���M0��i;�7uk��g'Tw��k�+ewliGX�����@�ۏ�O���O�i�r�j���ü$ewg����E1݆����.���5Ȫ�A')�k`̷��\o]��<��{{ڮ�o*eǝ��.�r��yN�)]���t�������;e��v(X�ݻ�t��:�Go/4���.���z}�S��G��bمpoG7�p]������R�Y%v�J=���r��N_$Tqk�y�Z�#z�#�lOQ�1Dk3�vZr���ѣ����]dp�]�&�ʦ�)�;z��	>�f�Շ��y��a��rDo�en��%�v�X}���WÜ�O�4���2n	�Z�.��^�q�=R�v���s��=���m@�o�ݭ�z��Y
�@��ָzD����yӑ7;M�=[378jY��w"�qF�Z�lu��΋;����Cs4ٹ���z�[|�E����Q����]���%�v�oD*�l5$��.��Ŷj��9��F�1�U�гcO,a�!=�ъb���VB�ҎL(�*Nr�چIMd7|�i�������]-!j�Rdak���m;ҭ��wl�X�k�躯aKr;8�vA'Z�W��������(EK�yٷ\�L3׍�\�)v��+�s���:Q�)�x4��{����e�r��r�Ʒj7{��n�����M«�\ip���7Bgs��p�z�k<�
���.�F+��8r�|hӬ��u�L�=R���+ͭu�0�tD��Ks�Q�۹I��T&P�ZȞ�LS]xhfa�Kva���{64I�Z��,W�`�2��ؕ�a�rhqh�(V�37M�QY�@U#4l�ѬYE��nU�h�Q����m+[��5��ڦh�jh�)t��m,�ط�E�:��ʢ"ɟ\N��A��[���٣�B� ��h�,�PQr�,��Yb�*��w��.�P�Hb��ಖ�uo+dp�1�A(
!�b�h���k]kn�A�f�j[�T���ݨ�l�Һ�Of�js����QyMTU���:�IR�_ZKN%a���):��m"_DO�*�ģ��P;[q:]�+,���A�8�RMd"�D5Q��ʚ�i�V��w�nܙ�s�9%��b.!�)��L;9���W��&���c�����!���	uG�"ǂ<9��:�=)��C�y���g8���srII��G�'��>��.'}�k�����qdA�Y����ǬE=|;������K��6��F?�r�q4�4�.��Zv�4C��$��mD&�;#ù�D�S�C�;i�d�o���|ﾻϜmL�������a9'�rh��P��pu|m{�Q�S_3�-�&?�Ja�Q��Ec�C�?ƒG����:a�����#�A��C���栟�rӕ���j�Ѽ�#gua�p#����@�l^�^�5��t�Y�:D}�W�}阙���nhUի��g��,�M��0��5SQG�,�ٜu��X$ܪ���3�m�o]ܣV�y�b	T^R�'�yU���"�f��:�6��;�dn,2.!QDҍū�x�t��|YP�B��"�4�%�úWrKW��b{�"�qÚx�.�#�j���}���&�鯘
��4����ܑ�j	"�x*�x�H8o������Q�!;��gM�Y��ù%"�$9�O6�B�މ��b��>ZM|��]���><9SC����i��[��<�ʇ��H���qJd9��C��6��s7�O��]�!��a!#�9G����Hc��9��"���cJ�}<Ł�I�q�$3�q_Q�9��$��$W'�"˃����ܛr��?|rI�aQ� �`�ܑݾ<z�S�p�ùE4i��?�z�}�}��w���f������,�ˢ��ɢO�9;C�8��ώDʜ`ē' ~-�H�9�9#��x�$��ݾ�燨y,�����8����=�笝��:cNL�]��&�I��u`��3���
k����m��4X�РЪ�;fe�w|��$�lҳm�:츙��Dc:��bX�y�:�a%to0Xy٪.ɪJp�y��F-:��B\���e������ ��k��D5	�1Ë�p5h�b.�U��g!�Ia�����!ɢ�r	 ��!�h����$�gF�]��|�@�J�	�0�Q���� ��$���ᒣ�߳�˩�x&�,�G ���C���栟P�R��t�&]�BIL�Y�� ��8�ˡ��g�'Q�DWݾ�og���BfI$�D�@�5� �.�T�Q�(G��9U�=#$�	2���q�Z4D�i�r�F�s6_��I�R�L��	$��e��aT��L8r$�"A�.�	�}-�2�h�B_"DG�C�`�;4%y9��q�/��OuQRܒ�<D+ƎI(�#<z�Ax92;9��w���G֙$���AB4D�|Au�˪+� �C����.jC��p꟏\}u.�I�mW[�]�CY�ʱ��߾�W��2�/0�O�|�l�|��O"�տZ�݂�~�41�C�Ĺ�mh-����K˛e_e�lu��4�)�\�t�U��{�P�m<^n3�8H݂݈CU�Z���^�d4ÅQ��D�>e���T��x�Ap>�ǨB���Ki�OX��>�h��ѝ��}����&I��!!m<a�R,Mh�=%�xӀ�K��zQ3>L�!$��8��$�A&Ab$@�<l�e�6}�+�w|r`I��^�!�*�$D|9�@�Zs�^}��E]y�|��$̓3%>N�q��BB4���/$�r9�;lϻ�ʪn��kL$̐	����4���ܪNQG�$�s|����[6&��9�d���&�8��"�hͥE�^ި�2@�	3y�'��
�R|Q�(C���NY'�߹�'��bd��c��� ����!�yQ�7�9��=>I���^8�Ȓ�@�8��W܃b=�u*:� �iꡃ��y�gQQ�r���>Q�$ag�]�W���b�<~�X�.��h�dh�B�,0�l���;ٖ��K'e
���rO��ŝ7-RP�Uf���{*���ٕ� ���qҋB��c�`�5���% צA!�YU��뉒eP���d�J��Q�^T�1�R䪉���	���9��4���NYnQT�D��
Jϳ�u�˾����o�eEav"F�$3�<l�#��7����.��ɟ� �&���)U�D9B �f�鈒m�t�q?RZ4D��I��@�0㙑�7�<�Fw{�ϸ�sQ�$�C�%@C40k���?i7w����x|HKDI�Iǈ,D���%j�0Gq��b,jC	7�xC�O�$Dp��@�Zre;x��N��<|}�OQ�a�C�F�A�d��&��P�	�������3M���zK-ʤ�a�HEv��er=T|�ZI���q^$�q$�8�IB(D�d#/��ڝ}�5S�$:�q��cSz��#�A5�����l�~&�r�j�2�K�]	��ԐA�`��p��l��n]�u]�j�_X�K�x{���$���e�W]nȳ��y�^�;<��0}�	�0@� �.����Q|К��u���h�␛�y�w���cp�/I�F9BM��(ҋG�U��w�w�}��	3"ϐ� ����C�|�*��1�4�=����ч�"O�|q�W�B�����bm�L� �8�s@i�U�,�(�\"HE��8���.6j����`�-&Hg8�X�3|a��~�Ȯfo�6�m�AH���(�(D	��!I��g?��D�N0Z(G�7I�9b�a��IH�/<"�]����\�"DA�
�-HI&�h����{�_����q� 1�@�Dy��"$�A�^�/��֤F��s-92���㇒�fW��Y֢�j���@�� >�>]ɼ�,�(��g��탱_K�{[�=��,P��A��n��n�56�:R��C��tr�b�!,�l˔�xjeii^.����3Bq�w9��� ���&���D�Y�Nk�Z�eў��^[��&)�t��xB,����rI� �G(D��i�^e�})n�fWY?�'�U'(��Đ�탚x�$�H>�wz*'"=(�OC8�Ǥ�"4�G�4����"���qE�9BM�(�F�P� �Ϳ���ǲ���4���C��PU'h��Ñ&��{�oK�|ʣI�A�+�DD�i��(s���{�b�#��N���ܢ�|"HE�99�F��ܒ����h��)L��x��,E��l ��I�����\��f_6��G���&�O54���Ǽ�yk��ޚh4�E��9���JE��M�f{S�M��~�����ô������_9Sԉ�Ҭ�"%�!���b�Rs|���*�kHҳ^�6��K r�a�aGŖ)��Il���eUWq�)�juW�t�g	�y�ˎʺ��.Ѝ��\a.�V�3i��')��W/�!��@��/���,��v�k �&  XQ��D�]p�(D@���!$�I���QƟ}�я�5�H�
�.������9�9"9�/�l�_�eLŞ1��NL�l$���BB0��6���L=���i� �r�H��4��|[��G�*��^�}�r�>,�B�s㍲KF���7��fffY�3�aR`��!Q�R�4�H9��}?}Q�q3^0F	���Z8D�x��9����ʁ�s�'��eRv�h����@��}��ٜ�����Y'�'�4DJs��P�k@a�sG���"��<f�|U/�I�!z�Ih��G|v�����yL���������ٚJ��L��'n�8xxRk�]C}�E���Ǜ��>	�`1�S,��X肖6��Y�]ukr�y�yZ�[ޣ.��(U\š�}������b�W,ɳ�U�꫖$�YA��"��-$M���l�.:��U@���d�¨�&^	���0��"��sH>��R,�����*g��� ��&��54��$�x�y����޿�Ͼ_}�#q9�Ye"��&�sd�ŔO�� ��0���5ڐ�G4��,D���Zz��Զ��w2��<"$�A�H�G�j9�4��{kN®��X�ϓ��a��(q�a�� ��4�k�ww><d�AB$M�4���nU'(�b���䃦|���8ì�ф��l��ȿ���ڪ�������HATlR�$�ÐP����5��^0�5�Q�Z>�A���<r�����7��wwy1�/����>���D�����r֩�#另q��J��������6�^��|׊�'mP���h����j�P� ��1�In@kyi�9feZ���m>��R^��=v���g"R}�ݏ���V��;�r�Bey$q2����vD�H���=�n�+�p�QU�>��cǫin�́7`A�8*���Q�%�i�b�e������g�|�A<`��8�AE�4�lr�ɳ�_��ò.���<T��DB,��%�	��9�[I%�q~4E�9���AH���<A�A��b��m<P��ji6ӄ��qG�b8.|g���wb���d.�Q�,�X�$�zJ" �H9���S^����Rm��$�Q'X�!a���9�~[�2"p�a�At9"!y� �Nk7ޢｱ�<ݽvZ��ǌB�F� ����PA���^��I5�w���4��Ia�H�AÆ"��ז��}G�5/.B��S'��OB.�q�3���w�cV�<m,N���X�ҳ���*Ĩ�X���][Tv4R+3��z���Q�YA��~�����ٯ����*�ʻ�-�?K;~L�|����pݿ{�Dg�\g��}a�q�}��V��
H�������>;���\R�Ul(�kٓ��Zt����f�gk}�oE#sϣ��xm�Wh��Բ�%��c��ޑw]?L���9�Nq�VS�|%���(�F4����s9ʵ�Ox�?K��^�ʋ�5E�{rl	�Wo	�^��[܆�/�H�F��U���B���1{��A6j�q���;����v��%��ޔ��jNb��.P*
]�[r�!V�*��Sݎ*�TNB��P��yKە�m��WNR������/9J�R��]�t�p��l��On���\�z�F�f`~l��/8�Y+o��������<�\&?Y�{@㗝ܩ�҆)�3<�k�����G�랼
9C&�8N�g,��=�4㩱xU����XΙGb^����*�>���}8P�ؕ
�y)Kp9p8{�9B�^��2s�m݄3��-�_*�ʆY��|��ٟ
t��D�k��RLƩ��Q���9�)�M�����W��s���o/72�2O�nvq� u�Y��\�wF�m�������^�$�_[m��˖�l�Iw����In�3��O2�m�A���A��Vӝ��Ä�-�,��%��__[d�K/om�I-���w��ܹd�IjId�I$��m��zx�]$}{��4h�C�$�( ��+��|��euƜ<�>�Lup��.���t���(e�"�;GY{��}�V7����Q�$t=F�(�����Ef�;�^�\�����tXު&��;nl`��s]��]��ܽ��K]��ܺu���nm�`�ª�y�mp�
l0�}�Z�B��UV;�q�N�6R������Ω��ꫡx5��^G���Ȑs�d����d�#.8�Uu��PO�r�T�5���U�������Y�V�n��ɘ�����}vgoN�sh�Ș)���hɺr�g��U��*A[�������m�F�'�b���\������rЁ��*��D���:�b��/�
��EghG��	�ö��$�&\R;9����ËFB�s�7�m>qZŧ�:b�8���ف��(�ZG��W9�#t�*��/
qlk,z�Qպ\q��y;���:}q���^C��V9q����S�MX��\�4�z�39H��9N=f��fH,-�|��Uae=��[[6>��ri�o����2��aꪧ�:�u)���	�r=;a�����Gws75����P�/'pR���JAW_*w��y�֣��e6��Fu��(�%й{Rj�%kU��uˮ�ҁL�^W2�_����T�hCt�U�|DKu^S�ԴL���j_�\U*�5�b������9��5`�.�vb��k���]�j�A��d.�o,
�=�`۶8�EHk8�.�YYl��ڲ�='o��œ�Ԓ�Z\��}�{]�J�V��J����.Փ�6�J�N2 �2�^5U�GW�)��H�f�E��v\�l�(藛y����D�J�؅�jԙ+BqCd���d=y���ƭ��n�&�u�Z�RĀ��we&5�fe�j�Ѣa�A虮�fs)�Q���u�j��	KiQ*��lA��޲�B�F9a�櫱X����CyS�T�O0��0�� P��s�B[�?h���{�B�y��CPۿT-l9��h{U00UC8�)���m��J1���n��m��F�7H�e@��%�!J��Ob`(�Gmԡ-���(p�c�9��#/�ō
}uwʹ��p��|�S{���]��J�-�ҙ!�ͷW6���d�;y`��xD����������T|I��LH6ܧ�x��ò0�L��F�L3�|l�"�p}U�B�z�}��X�a�t��Ta��!��x㙰�	���ھ���f�K��� �"�.�(DxqHaZ����|L�f0��k(�%�|q�W��-��꫿0b�M�枓�9V9ER�G3_�rs��3��}`q�Ñ#�cY�H��$�h9��]��]��Hf��x���
E�EaD9B Ҋ+��/���Nli3S���I�"�Iq����~$�=�%�wh*9&�,C�%�a�
�-I��o��HۅU4�H�QgX�!x��m�c���q�����٫�k��!�Jگ�߾uK�>{�Ґ�;g�> i�!>r�*�^X�jV�oi3jR^��<c���*��un�T��Ī��nd8��}u|�@�r�>����3C��AB�q�[�r	�&L�Jaܭ��^��R���OE.鴠H�NT�m�Qb�OC����ĸy�k���",s�s-92'ox����[�>�Q�ux���8�AYd��NA�(G3\���oz�������Ko��YnU'(�B(C�3}X+�S̼`#�:�-I0�9��(E��B�7*N�����'ʾ$�9BM�+����Ҷ���[����i��0�#H*�(DX��Z��P�Nb�]���o�w�9b3L ��b�0DJ�9���e��wp��Ml�'X�X�K�B(��q���[��wv5?�0��F$3�$�h,��9�ޜ����1.�Q&��R,�+
 ��o���?Vh��:g����b����*�P��}d3�k�بj��-�x-JV��\�-K��Wz:�z,��VR=Ͱ�X�4p�(0�B���E�ݥ�\���6ݷ¹5u3V�s�vN����AwvΑ�i��n�K�҂�YX�l7[wV����1 ��0��(h(d����O��lGP]
>wl^V7$2L0c�	5����$!����E����F>f��a��Y��(D����M��$��3�w��V����?���D"d+>>��\"$�A�pm_�:���`�O#��m�&S�Ĝxy
9���'��s|����	� ��i� ��"m4�m����g{f򲡁H_[�I�(�I!!�>7l������ި.�j����>w�$�"�B�`4c��Y2�޴�|Q�r�8�OV�E�A(F�sq���h�k-�R�TJ(M��5������qw�N���� ����(C�I�P��&6:��_�������x�%����������/Y���f/O�|[���o*�4�h��&CD0�cE�a��4m�:&�ѷf>��7��G�V�G����t��%D�.��7U�޽Cb˥1�g��X���^���O�юϠ�9zY��1�I��:��4MC׉9����2�*�(�Z"HE9�y����"��[7�x���#��I��H�3�A�������.'}�]y� ��>3J �(D	�|y���N��=_{�R��t-��-"HC��v�-&�4C�����mD&o�C���0�M��$�H$��9���~��|߾�Ϝl4�2�2��<"$�A�(�������l�f'�y���'&S��>8y
qi�����:�$$�]$��&��r�H��C�>-�`����y%�U�����(,���!�Ü{l�т9��~0�v��Ȝ�	 HI��q�>��(D4�F�U*�%(/��#�<�)�NӺ���ݳ}4�#H�)����%D}������̀�;7��Jr<�,�����{|�� ���EH$�BhK�hZ4�$�T2l�p�,��;xz�Œ��i|o5=�T/�c�N����OtT=�U�L�)ηWaӻ��B�@�cEUI�.T�?Qt��iS��d�T	i���}t	ĽE��5��I�L@�Y��Ԩ�|"	B<A��'�O�yoL�!2E��G�G�J(M�'�\�"h��x�u���O�	 J�� �Û��(C�l"��a�s��|U}ф��Rdɗ�9��YT�D�� r8s� �NY��}���I���4�(,��_}� �YZƿ{���J�3�x����A~o�<��anKqGo��N������3i������-&�>礡��g���8�&qd
�mHI'�q�,D���p����d�����<"$�A�(����jg9�~F���뻪�����v�L<<�8�4��d��Kg�����U�޲b>��|���L��bk��:o����*�uTF#�<]�Z�rI^��v��	�8hѣF�0�Ŧ)&Χ���P��Z��i�sx�d�^��y�}wj��	�肹5�70˻��N+`C��R'����nTj���k��y@�q�D��R�q&x�K�:�H#l�B.��ݡI�C6��˩�0x�ϥ� �"D�|���ܪNQ�q��L�3Y����mþ�KF�]�4���dWݾ�m�fVI��ZB
���QXAG�r�p3Ͼ��UW�,��6�qz*-"	B4��9B� �+��$�)@&���a'�(D��ic�����4[TVh��i!q&AB M�9�����8�ogj��T37�>��$�Q���,�19;9��Wy��DPw�I����Z,�+� �5����dDm�Wk�	��榓ŸI-�(�,G3Q6o}��ϳ+�#����E��M��B$D4�I�����1�mn�i�k �p���?"۲?"
?z���{µ=�o���D�$�!(q��$Ͻi��\�z�;�����i]��U�������.���Vܝ��m�c�v����Z]��-=�u��i������M!��.���؅+�`�U)ݴ�l<vڣ���t�W��*�TQ�t"�T��KM�[Ip���#��i�Z��M ���H���_�"r]��a�L�|!�-H�xs�s-9���v��u�}�;3G�Z�<`�8�4���/$�r7���(ϻ������K�5�%��T���,ts�w���1�!��8βKG�$�q�=%�͉����~t�n�)�RL�QM�I?A(�� ��r�8�4�53a�e�?G��ĆI!!�	��7xsQB$�#�[�"�� ���}��L����$�BI$!$�&��UZX�����ǡ7X���@�8����)6��o��뫟����ZB��V�Z*֊KV�ie'�t�~�P�c9��6�*�(�Z"H�e%_������}�}�|�I&L!&d�I�&e��j�Z��ێ�q���O�wz������ik��=tߟ�ze׵�����`Y�8a���S�G8GڽX�.�S`|B	^l&��>G~��r��{�f�p�l0Ŏ���!���ݭ��X��ѵoXIeivޖ�WsY]�*��&�G�
���]��/g�ǳE\M%���{�TYH�A;6k*�V4�:TE�"߄L��)T)$y�R*�@D�I �vj*�HS^`��k|�-ؒJ�-]�틩��~��L�4IU[{q��^�;�㧓�Q_AP�]�ԺN������K|�i�K|Q�E��������y�������q��4I��.J" ����Rs�G�������G �N=��2le��8b�>�u*"F�<!ωG������NL�oQ�����OyS�p�$#� ����NA����\q{�w�v]�!��<���ܔQFx��B�<}��x�QC1��:�Ih�4��x��"�9��g1�>�]�c���/�#J����!��x�K(�p�^��n%�}��|��qg�E�H�(���c������k;t~d��Wu�Kkz����oy@�U���_A,��������|v�Z�2�P�;��3�ƈ6�%�@��s�L�n��Ɨf�[v�ӮQ%V�s�ŵM`��s�vͭ-D��{k���oQ���-��;sj	h7�0|�B˧�C!D ���d_!t	T�K� �,�zߠ��8�TB�A���X�HK�V�/3	H�1z��K �� �]�����{��a�X�bres�OAֆ"~ߥJw���D�8��.�.�(�\"HEB�G���5U��m�tA����H��x�$�o�0����d�U��8��E�EI��6�5���>�}����$�����b,D�㏇�e����/��Gu��k�9rP��*l�!$�i�y���=�3�a�QX�!i�V��D�!�<�f*��/�㺡�,��Q�M֜�N�|Q��+O�D��0||"� ���r$����&�7ɛ>4�2�?;�fd��I�(�����4�тw��Z���a�^ž�@Sw��Ͼ%J�|C��wv*Dj$� 3��%����=�����v��b���1���)�2�$�B�B���t�uU��v���kKZ�dZ;��AF1ɖF��坻�:��v�ʑ|�$EL����H7�2��ںg���!��Q��v�5�Lzu>!U/lG
�	��I�.�p�̊�Ȉ��<�|zJB���G��s�xDs� ⳏ((C����(�NJ���m�/v�=�]N5L9��Q還�xEɣe��uiV����8�Q�X�92��OIB9�����&��KQ�#����r�r����!@�#��q�修�\�x񸜉��'��@��V�9���Ͻ�B��32���G����@�<��an��#��Z�<;�A��qh�C�>�,�X�$�o}�tLt�E T�jBI���I�Tq��otc�M��H�
�.��<"$�A�(������:;����L��u��;����kד��i�T�k��Ϊ́b�Ά�Vq=�r�c�P�9�0�`מt�Mozx���
���,g}���ޙs��t��[U��aɧ�5;�w��&��;}����%�꽽����{�͝׸���*�S��&�r����n�K�!p_7�jR���׏35n�y�������a�w��t����{�,��[->��3��m�����R�)^_Q��1��C
�6�q"ܿ<���{;,ee�0�����M!��K�\Rl5��t�U���GR6H�K�k�
�:�쏛bU�o�����3+d\p$�%��*_[�)��'~T�s���Q����Y�vk�+T˛�t��Ǝ�]*Ld��Q���	���x���P4ϒ��ʭ��������9w��u���ę����,&u�-����7�y�(���wzS[R��� ��;	~Zk��!�{Q���>��C�%�Ki}������_L�-#-��W�P�u��u!#2L�f{�<l�����"��(I,z���^K�7P�,�,����|��[�R[�BvZ��J�*�7
��;�Hl�H���:9��)X����!ܤ��f�`��_VS.�Z�I�鱐�\ދoo��v޽�����y�}��� <tuӜ����t��˗.I$c����݋F�$J]�]�'0�	$�Ir��$��m��$��n��\�]I$�]���嘗��I$����˖�l�.[m�K�^^Yd�I/n^�l�I$��m�I$�Is33�:���;���Io3<ݚ�I$�wd���7 ؜��[٧4D\��M���lɹ���n�.�ZlQ��z*e:r�Y�=�[�����|�M혪�w6#���E9WhC���8z�e;y)o��洇Ls�Mʏj�sfM3�*n�.���{��sl;/�r�w,�7����/�*p�ޮ�72�u�ۍs���7jG��9��q�s�B�.�r��Ju�F��G��Tm����Nc������������ǲ����:V5}>i�*����X�U�K�W>/T;��;��ڤ*��:���T��QG�I���cݷ4[�zVǲ�攼�
�{��r�
����J7&�)1���s���wĎj��f��M4���A�9:���W�Ӵt�Xn|�5�U�F�u�_c�������j��/C�hj���D�qf=�ݫ�GLaJP�1O':R�y�ܪ�WHgk� ��Ӿ}LKO��RN�uͧ6�r#'�
r����v: �:$f��E7b�c*�}|R�ʓr+.��<�w:��t�]��e�*GMY��0�S�bg[L��r\�V��Ӆ3vdrXݐZ�wt��_ت��f�P�s/iL��O�2m���H1��X#�d���E*oi�c��#s%z᲋�7e<0]���\b<��[�TȜ�j��h����Ne�֥�&��y�w9C�ڻg!�ϪЅ<X�+h;1��m��䆯E�J��+�ď�]�
q����|���Eӂ�E�Z����wP��!F0�X����k^�ąVĪ�)iͺ�fQ��Hn�v�4h�V���*�^�z�Z[A`�$☷���t(�R�"juG'Dޝ�Z�.[��bŝ��uaq�� ��w�+D��.{��G�O-�r�,�wi�X��A=�si1d��JǭDb�y6����kH)l��i��G�Vvi�1U �)��Q�`�Q+RK]br�^�����4��I�ε�"��C+vQڼ��W���*�B���S��)�A���	I��i�uH�cw��]�׋��\ס��]eLB�=[4����:MS�9�f;FV,��cv2����ѡp���ŋ��{�f-�wW]{'[�x��ѷ�˜{n��۔���vv5�@ث�<%�T��b�ikbτ��>P�<�r���� ��MQ�����w=g�b����=�C$�d3g̊�����4��}��2�a����zӓ)�(�(q�a��m�v@�c����* �
"n<�I�nk]�o���U���G�P�����-&�c��w��{333ϐ�,�
3�eA(��ҍ{���򸙯#�|q��d���x��9��V�+e�ꡛOC�@����(M��rP��x�����E��fQ�`��res�OAB M������T�3G>*��$�P�#�<Ybs�����2��c9�u��- ����YZ͑��^"TN��a�� Mg���L-�$GiF���^>�����{A��@��{�-��<~��:E^y%����Q�k{OH����A�9$Bǆ|/��Cfc�Զ��5�E1�=���k�{�V덅��oif���˧ٺ�E�4�J[�[S�A��(	H��Q�����$V�$�Gα��|���pQ��$�QL�J>�Y���x�_�T3+����m���G#��}e�D�!͒�pQ>ߠ��19�'*k�!$�A�GAb L�f+O^}��]�$�Ì��:�(C�|�$r<9�L�a�n��Z_S�]q_/��MFxR8�0�m�Z9��M=���=�$rܡ8�4'Ź(���q����<�D:,C�q}d��I(Gz�O��ۻj*���L@��1����%VQ�9B8���S��^y�Mgt���$$�#H(�"�8
�o�<D�1�'�,�ABn$����@�8�,s���G�\��3��)A���B�K��@��lr�e���ayp�1��Yɵ3(NjK�?ùH�?�P���:8|~�@'�>��)�^��r��,�΃�4P���@��Ō��l�M�l��'{����ƺ���n��E;���R[%��.;�׸��͙U	�x�� �+:Ǖ���}E�k�4!�,�ŤϬ�l����6l��6���dS��P��4媲w]Ӝ�L~?� �	����B(DdYbr$vsN[��_;�jdɒ���"H����*��D�A��b���H�	���E	�(���Kp��Gy#����݊�j���fHt8�W���bh�9�(D��M �}E5��{����I	�ݶT��Q}��2z
�����#�j���3	C2V��4C�Z(���皙̵k7޲����=��g2@��	��ŊB�F�}� �aSA#���7�t�^��Ͽ�M�ڲ���'�9�=�ܔQGx����V��̼�$�ZZEl�*��7�o�~=?��J�GPP�1�{�]�R�3<$�d!$�&L��	g �2	E�|�~���-�^���b݃qZ�c���D��{Ґ�ᴂ�f���B|� \ԟ1�oﭗyl1Ns}v�|�]�������1���In�}Z�ͼN[G12w�k�bM�r�ƥz��λW�uױ^P{KB��D��ҒD��9�����UK���Qj�0�s��nMĒ#$N�z@Z��P`�U���U����0@�IL�ύ=A$�AE�B �@��z����x��6�QJw>��G�(D��<X�bs�CL���/U]����6!q��B MËOI����h�#����N{�&r�ﯙ�&I�<#�I�Y�r$vsI4�b�]��]ŗK�$��Y��*�PZ,�+
 �(D	�(���K���Ĝ��a�"8��E����O}Ò컽q2%r9ȑ4Ib�(D�� T�jNc�sm���V�EUk�G ��:d/z
�p`�f���Υ������$q��is-D&��)8�߱�u�غ���d�G� ��G�MB�o��2�P��d{�^k���6�w���Zk��<E8jiޝ�fٕ/<_�!��6D��A*:��W�nc�0���BO��T͎��/(�V֞���vv5r�k���f.�Wf=���gU���֩Ok(������)�c|�:�oUᵸ��R�1��F��R5�JzDM�R%Ek���ђ=��6���E|���`a��Fx��B������S̼|��q=��c�$�z��A(3��j~n���	BLY�yW�`��&Ï"�1I�u��=�Z���}\æ��x�(Dd>�F�&ӆ.���{�{��d �>�@�8�9���B�M�����Kϱ1)��qI�e�]�QT�$"�y�N<}��u�����1��A�A�����&�Ab$�1qNx����2L2BL�C���b,�+
 �(D	�<sSI�;�I3lԁ!���Hp��aĖc�"C��Q�Z8h�Tc�n��~Jʖ���8���zN�.��02 \�3�5W�'���z�[��?
m��H	��ĵ!��J��W�� ���4��ې�E$���}:���7��|L�I��(��9�����ks�"_ea��#�U�Sˬlv��ݤ���ʄ]b�wj�F�a��J���ǼM��r@�����j�E�6m�	�#��A�ߜVq�H"-�م�ϭ�3		K��2de��(�A�8>��Ft�7J���$�ZX�$���r$v��
B�&�������h���q|A7��*h$s� $q�M8p�g�{튺�Ԑ�y.	)�Eqf�:(C�|n�'&o�3�{��Mx�$$&�N�!Q�">�򍒑L1��0�|�d$*�����a��+���t��ݧUe���Np�#�?�Qu	���&�����Z�.�#)�d�G�QF�Yc��ɔ!�$�
9���ؒ&q�D�8��/×c�U.$"�A �x�>��O��}�ȑ��0�
dXA��	�>���7�Ux5�Q�| �{Ƚ�˱g��~	W����Ř;Z=�B��{&5�Nֆ�<4h�>�҅c�I(cJ�D��\q����bS�%VM��39���8-�;�U��grw�<dƕ�j{R9,��a�0���rh�P�U�Wx�0Wm1b���&�}�(���C�"�<y����8o����J��3���a&刂���6�E��V�sd�N3R�x���*l�$"G��:�}�������C�&B������Q4��9"8��6��(��Ѩ�y���r$v��G
B�FA�����T����9SA�D�;|kA���0|w���$���!�,������=�I�;v�wm���ɪ�4�#O��A���l��+�h�����3�$H���qgH�����x�O9�ͧз_�>o �G� z���
|I�%�w��
i�����ۑf~Z3���=� ϑ�)�L���&�*9b�t��"��>�;"z��;qo��r���A1���%��3v3oj��8G��}m���������g�YK+dV�RJ��\�%��u"i�R��%�g�R��_*����ۍ�ٗ)�!�3Q�^�����<9Z��B�M��m\<�����lf?��%�A衣0�!E�8�� �Ns�Y���"0��AƙAb ��� �Y\?�{���>���=���&���M&�#M$�����߰����_@�G�C�E�e�L��9�(F�}���"eM���,�Nڒ#�A���@�=����}�����4E@�>���i�����0�gt�E��VrBYI̱��(�(q�a�� �࣏��R��$�]�g�	v���>-�Eq��i�F�9�2d`���s��0�bIB4��}�#�����o��?u|�ꋬ=��T(�<C�����<ͪG�k�?H�-�y].��BA�#�@B�A
u��W��O:�g2�Ӯ�]S���G���c۵ױUvI�S�Ns�&�mL�Bs�wj�v/]�im�s�fUU�x[I|TfR�h��Z�\�QUTͻ������}~���d�!!�Q��@�E�H�������g�}�Ȫ�]ʏ	$&�N.E�␒P� ��P�#H �1�|�Lt$��x����I�.J ��X�1������P�3�����8� (���ņ����8����o��c�/���$"�A ���3�#��4�m=S�x� ��- ���e9Ep���I�{1�6�k�0M��M'Ź��>$���1��q�y��뛞�N8�nYe���U&F�B$C�x�N����ޔL�����RB$w4��@�js�/�Y.��3 6���DC�!�s��0e�#������0��~9�@�Ń���5ȱw���������\�q�YʸzUIT9Dt0ƍp0�p_ �A80��5�s��Ur�푔����7��7.��Nʶ4k��1Y���7�1�'S׷-��5q2L7"j���˲o��&]ӎ%C�ř7����_�y�iI��)
q> ��Ax9SDszQ1�Y�wASO�3 �㴔@�L-�Eag:8o�������F2,�:�>1ؒP�(�ѫ�����}���,��p�JE��!��q���YF��?F'����$�#�	<����(���a3�DG�Ţ�x�!DA��X�bs��7�=Q0�g��q�4�
 v����5��$|�� 绿~{�i���4&B0E�Yd��ȑ��(����D����Jk�XA]d�)�+�ǂ�@��f����+E�4�c����K<刂q��0��G���X����M�ʽ�z��O��^�(\���}���)�����n��4N�)ƊwRf��۴sU�#��*��-�/h��;�鯞>�p2�4�;�r�.��H��������Wifp/.�LÒ��fS����xyl�0;���tck��uX��əZٳ~qV��Ȼ�Y�z��9l��I�o?-�0���G&����S����9�F����S��s�г�'m^Ֆs���(���<�z�������N�.����Tج�ݓ�Xx�=�/��	2��7�y������|iU���o��~�����9��6��U\,�a&��~x�V쁎���(w���^v���5M9�6r���]b��7ŵ=��Fӣs{!�'�ۜ,���wf�GW^t����s��m"ϫa�[Qsˡ�ҵ�ۻhl*}%rȖ�Y�w���t���U��s}y� ��7�"�+��^ڻ7vޮ�勒�򞽞 �̣�����[L��E��V
T:���YBHk���Y
����{��t���o4�ޕV�5^qE�ڎ���
�Vo7J��`]�݋�����7�����tuۃE�qjU�$�^�[K��B��	 �x���$���N���Y������e�r��˒I$��}}l�r�m�O�yyyy$�[���u{y�Ym���`�� ��LM����� B`�,�I/����l�L����$��������$�����I$� �p������W�kvN�a$��R�%U��MV�F6�9nf¹���z����Ȋ},9��}��l{Qn�О�U+/w�=#�ܭ�z�)ֹ%V'ٔ4=��j��)������e>�*��hӻ1vI�����B�N(j�=�gv�ݱ�fM��ˠ�?�G����Ua�(��=��Wi�綫v�={�P�T���.�.mb�N���镎7w��*���q�]R�'M_n24�6�@�ʐ���J�}��6H��}�Y�N��Qj;�{��׋f\�r��ˠQb��{7 ��NI���]�p(�ϝ`�ڨ��NVh������s�T�C͔"��B�V�w�ō�]�T���{}z�<��#�Mǽ*�|�)u�-J6uԻ8�9}�)د5vǝPJ��e3z���]�7$�^t�U��F�V�d��)�oOb�J��Ol��>ĩU�;��{��8���j��g,�	�{�{�����N��i����e�j6v��<JF9��c��������$�]X��
_��^����^ujO+�^s��2�UZ/����k���)m<�.�g^i�-���q)�T��>7�hH�U��\L���ت��zp�@^�&�*�F:�6��=ySH�Z[����vm۩��ñi���O�����i��d��y�d�Zm�T`ǖI�$�nf�ZrL��˘y�r!.�^�'[�OAdf�V|����5N�勫��B�X!�s�=ɘLx�a��%�7��X�[����i�e���8WȾ�Y�R4�{L�]�?wm��`�!���a�m�8����4R�i�扏.$!l&1l����Cu����2VZwc|�.���\X�Vʘ��2P���f;Y�p�`�g��G.@�Fk�5wZ��c�,� �qC����0��k�v&0�mc�R��>P�Ҵ����ᘷTS��B�U�D8�2� ]G�����*�l�0e�BRW\�S��$�IV��ܝ��E�h��/B��%R���^�U��K��w
�ܛ�2���8��]sf��vn��c�dفA_1]��ʵP�E7o;S���[r�ʳ�u�֧�����F%<�X͏on�=h�#�A�U8��FZ4�����=0[e[ۙ���V4f��81���	��gh3�"����SY��k��`�)Y��w�촩�	��],��$�� ~�C� ~c0����H� ��"��'�;�����5�b<��܃�=%��2l��1�88�qԨ��r�9"�8Ƙ6ӑ#��(�I�Ox��ʞ�܉ qY]�_�*h�z�x�;x����;x��,�)Q��(tP�dp��C�J����O;J�GPP� ��9���<��~�i�b4�>(�ABM��6Efb���3g��m����F�2�,]/AG�	��Ӌ���ȏ'�6C�A�ac��ɔ8�Ǩ����rQ.�m�$v�ťIv9v9ER�B(G���r��w��Fs�[�fHK�������d��X��J���;9*9{���܁B��y���4]��a�1�wF�ӽ�;����s��O�t|kV�虷:i�P�\�(��r��Sf]��hqw���p�j����wL�ba�^�AH�,J�[ń[�:�H�����5U�)�>>0�؜����Ab �������z�Ȯ��a���-	�g4�p��/e�D͒y�GÜa%�刂����ѭy��R�#���Fbd\�"D9�)�RB$} �
���o����|ϼ.$D	���`��a�Q4�ls����������(��N]�&Gm>(�HQ���Ϣbg��qv_Õ49�@H㷍 �k�O��_�.�ә�=0��Ȣ��<P��9���8f���ח���cO!z��A� |��R4���y �Ox�9BMg"�1HI(GF��c6��2��l��0B�T��O(5��|}���xW#���>g�}�ڇ}��A��e�K:���F��
�b����܇�U5
��_Mx��Z��u�rU+���܃[��TS%�U]qs�[��%k�G���	�e��ʈ��nZ���r����B����Rr`��p�ي�T��0!����C��� �!��E���&����#�IdX�92�9��������eUP��v��GI�9v9ER�D��q��e��d��]�����ȑ��Q�XA��3]l}���\�wś�j�"�a��$�܄s�<|o���s�|刂����E�iT�'3I��Qӆ��aE�)smD?�Q�5���O����1�&���&E\�X�r��DX��/�l�y�FO�� �S�iɑ�(�(q�a��~��&���禂>�D8���O�r���nl�m��Kă�:j"C>��CJ6���>��
����t�=U�*gXw�sH���Don��f�y$B��}�0��.v�9�6��ݼ��u�6�U���y������[�X�o�֗�[�����0��1��8ⶤ
���$)"�-�

���ܧXK�[//��cŔ:(C��>7l�v9�>//ݽ�t�I�a���cE���Q��8Ƚ'�3�b,M�}"�qHI(G�s��z=[��������?�Q�	���.B��Y����n�"�o�x������QC��8��8h��qO�G��ϊ���!"���A���~(}3g�s�0�ZA�Y���`��G���⨩��>>B�g$��$�܄H�If�5����N���!jX��ݏI��,F��Q>����qω8�]˵0H�A�GAbh"�ڳ��U1]s�5
�K���IZ����	���T�WL:�G�?���r���E�R���A�80�A�WB��(;��J����ʚ�Y��**�壻Jt��r�]Q2��ؑ�
���u���fv�4���:��%��PB�% !Q�D�/�I�%摗� �WU«��52���6ß�@�=c�!�����l4��}���*n�1q��|Q�HP��H=�Ax9�YF���޼]�!Ň-��ܤQG�`�W\I%��y�q�b�s��$��%�Q�I�3��ow���}��Ð=Q���+(�1�Yޘ����õ�Q�/��HI(F�z�(C��s5Y��"c����o��7xE�Q�q�X�F��Z��}����]$��it@P�,=%jr���_޼;�˺�4���i"��>8s19h�9��6�Iy���c���* ��CE�k�W�y�U_�H�Bt�H��:Ǩ����{t}�C�@��
(i��pJ3�f˺$5����ņ���r�5
Ĥ���Cn��vq��UMͪMF�+��H.u���*X5�a��'R���P�Ffmٕ��8�TA�dM/# R
;6Sq�<�<�l�תbX�H�LTd�NT�,�=�e�������E��h2 CF�Y�,Gr���]�ت��Nq���W�E�aT���H� �I'��׾�AS�>g��Pc�X>`��:c�1��#�j�7��"���x�ħ2ӓ�}�&���{���>i���8�> ��Ax9SA���7�t��w~A"PY�4�)QŞ(tp�Z�w�����mò�4�bIB>(�
���[�/uD�f_���H�:d��+(�NP�a㍓���(���?w�qu|�|o����QP�r<A�o1���&_T�	���zB���<X�b����k��E���^�g����F�2􏁺c�.{i{>�Ǭ����H��S'H��Jd��MU��>Ԥ/ٗ~B� �|<�`1B���-n��6��IkT�EQ��6�Jzy��u����C��T&����uԑ-�=��ZHU����> �~d��(��E$�M�
�>��!�Gܙ���/U�;t)]U�3l�X@P㶎-=%y9v9F�i�~�h���g+^��<#Ǡ�M0sq9h�9��m~��겮��c�Y��/� �ܬ�Ь��6��Q]�%�[IĜ�%�r#�|Ig9b"C�o�ğG�䷾���S��%ز�22K"�$�s-s�O��*N�>f�@�Ae���L�zM��1�1��/E
���H�r,��Ne�&Gm$�A�^�y�������G� ���r��=D0\��ݝO�W|xG���)Q��(t	�s�y�gz�d�n#���v$�#�PP� ��*��{cf��J��\E����WP$%���}�AcoNZ���%.{!�z��%�w�G��˽a��6�/s�J ��P�����X�c3�oz�-q�
U��6���9����I��`���k)i�����^-<et�����%Yoi_�����[�yz�Ӿ����jԔ�)�J��(�q$EZ�]��T�4S�&�(F5�qQGߏ�&|AF	��l<x���O�u���}��{ՙ��GB<A~�E�@�PP�N�W{쫧��4���A$����q�6�9��O�/lDd!�8��+��(��MC���	8��k�מ����i&f'-'<iF�X� G0\S�>/��|C�ɤ�dc���Z�&s�����܈�H�����9gY�"!$9�9\��9��U���>n+�ȹ4D�r��%��S��9����׷��ﳽ��x�4M�4l��	@��C����׬:��>#�,���rdv��
B�F�ߖ��IC�����
��B�Z?����3����"%!����E��46��c�\�X���8A�5wd�(�� 1Ч���x�;�f�X]�͹�H����I�ѵwTV<ڵoEf��p����{,2!�dYd=BCG�>��h���4�K����m@��:[(z	� m(}V���.����y�h���ʚ��	��H9�p�Wl��E�]�,r�r�EY��탟�I�q���{��5&�wb�B>2�
�@�F�H�c�ĜY2����A'	��m>8���$"A� �`�'��.���	�� ���X@���?����������Ǉ(��$����q�6�
8b��ؒf�"nZL����8�MC��A�N7�>0η�7O�"q9��s�(��� �Y3}����]7U� (�#ß�d	����)0�%��={�R��~<Y�a�X���s��Z��cJ���;�a���V}y�Ta�4�\t�m�<�F���
�{��J ;�i%L�c��iW�m%3S�+1�Aha�0��0��.&�V	�b����L�N�����ֺwE ��ܳv�2�I�uf��M	x���ER�bYV�aʴ�(�@��Q(xd\����ȳ�0���!g�QG�o�[鸽�E���4A,���a���9�$�s-L;�>(�8��vzo����>�f���D���I��x�(�A��H�f�8���҉�� �|��ϓ�#��p�(C�A�19�T�Oct�z�.h�u&s��|[�1��_}��]U��1IF�(tP�dx��ec����W�ݷϓy�|���g�
�9����E9���-�z%L�30�#�5�a�+>�$"A�z�4i���[��H��AG�	�<P\�9���q���v��x���(Ej�%��D�;h��d�>��&s�ə�������,��4�c�����A|*�V�(����-�'
"��Ļ��%�X���r�o��<�����I��B�/#���^����sC�罫sz�4�Q9%�g��K�;1VJ�F�̃%Vo�#��C#U�����޺;x=�'{2wG�7��(��e�w�o"���M��O�6�E���u堳��Rs�����9]+��D�[#;��
��}��4�^��ַ��F�*�ݢ�A<���=��>�g.nñCb6LJT-c���uv�V�
H�����nP����f��[~�y�̩�gl��[��.�T[ծCN
��?m�uu߰���^>�{S_cZe�D���"Xb�-��{��{�}�ޏ����
��	��u��/&צm���o��wfԇ��
�n�膪�зj��cRQ�q�U[A-u���T�ˠ�{�*,8k{��8����l�vn�Q�4���`�Lܭ��建�C���|o�QJWf��T����@q��%�U��gJ׃U��g��З-%E�ǥо��֥y�2}X�Fk=$���޷�����F��z��\�xюT��RQp��r�Bm�����Kė�&�ƾs�lC�.����#�Rq���GyWx<k����{ΰ-��N���i�	PK��N��W�VΟ�;��Ӿ��d�T�J�z�8Jͧq�m���9%��$�L�.bI$���������xu��}�n��>z4hѡA1�6N�Z41$̺�<�������I$�I/oom�I$��m�I$��W9���^^I$��I?9f%��I$�w�r��%�[m��o���Y$�I{r��d�I%��m��$�I?�˻7��� ��l��RI%���o/7�uH��2�ZfX����D$��b�5��7L�Ht[9Q�?7\��e]T���ݡ�1]���W',�L���k4[�*�P���(M�r6%&+"r�w�'�����-O{U,�WI�"�eQ��c�H���xs��Jq�֕v�E@���7u���)}�oHn�'BJ��jS����mJ��˓���m[�o����{5kj�zm��M"Ҟ*�v���kŽ� �U���{�1n�բԩOq�o��:1�]h)ކ9�r<�n�Krj�Y��K�YP�f挝�²�:�a��jB��C���]u5[suk�wH��c��x�ntFj̸��������KD�Yl7{�X8�D���]��m��L�nf7j����yZ���ħ��9"��n��4g%%-��I��r��*�UjM�I�z 0���K^E�p����'�WEkgv��-���:�IL\8���BRob��{�=������3�������^�4L����t�S�؋��=�m�i��&ԩ�m`�)s�֛��ͫ0WR��N�H��V}����α]��=�*�2�l�7��Nk��ِCA�ms��N��sf���o����+ï> m�OL�D(�6���e��o����8�tq�/c�HUU1��:;�l�o��H�H����y��4���3��~�6FA�S��G�i�y�GU���in(�f����
!G-�ھ˲��-1�0���w ��ض� ��2�^�m$�����"Aol�v�o�4uҽ�P�D�nI�S[B�uo]s�TlB���Z��/b��V�}��{I�� ʖ):[J
�*<���N�z�F��N6�(MK���T�}�k!��$��T��dRR)�V�-ǕV^�4, [�<�ڪݩ�U�
�jS�f�R�7Hml�.�xm��:�%J�'«�������.���[��&�,�n���J01O3v6���YO1}�Ȏ��ȢY�"�el��0��s�u��KAu�Av4Պ�w�P�"­���j��՛P���G	�}]j7]��U�of���/���q,�1LB!U��I+51[.�
A�q7y��=CX� ����
%QɷuO(9��ΰ�v�	����2v�{�//R�'N;9�˵�7C{��,З�w��[t�i
)-�S:P%� A�$���H4����D�n�nI�Z��L4�x{���r4����7l��r�� ���[)g}�}�����_�9g���nJ$sM$��fzww�32����fa��I�(�+�e�I��,F�}���"$�f$Fqd��m��Gs�=%��L�4����\�w��g 6��s��Q4�,rD9x�*`ߑ�gtn�T��)ˡڋ(�(C�A�d��}�}��a��a]!��!"g8�qzO�r�Es7q��L�x F:<!�a�YF�I(F���f2N.�}���̮f�M�����E9�

�����9>���M��8��� �mP�!� Ͻ�}�..��W��q��|�!wQ�Iʛw�q����}�	U}9�P�c�e�]P�ˬA�A �a�Ƌ�o_M�Ό��EW'N�����o9���6ը�c�J�\��=��PZ��Ǔ��U`���>!��=z�]N�T�O:1�D��C��t�԰���/���CE�&�J��@� �#������뻳�`_'>�q�.�
v�qa�Q�(�8c�8�{r��4!1����?�">8�br�H�9��͸P���Ĝ��	�
� �ܮ�Ь�F>���z����`�H>>"G��%9�Ės�#�Yg~~���白I!�5��e�U&F�b$C�x�I�>�:=�L��7�X�	H0���4	����ls���Ed����F�E�X�$A�O�Ne�'@��>������>��"i>>,R!���z�/*h sx%��3y�EK�	|&rJ[&�"�0���+�K�Mm��_�E���d�(�'�l��^�	������z�p;$X>>�J��k�5���ݛ��*t�A�*zUVb7nf�W�t�*��F�Z���,t���!ȳ2��Ln�fi�{���e	ts�n��G�/أ�*E"|	d#�"��CL�
/�Q�1����^f3p�?{��/���d��&�sOIb(GWi�s���w�:ae�@��R(��<[9BM�i�pQF��ttO���JD��z�(C�� ��7�9��=3y"D�Q��P�x��3�<���ǫҢ�����w�3�x�J5�-�4�M#�������ט���ň$�(���'-4�i⍰�g�e�3�b2R��Ae�_YhV@@���l��N�����(�L�Q#�Ig��	!�9�f���y�����6ʃe���ȹ,D�rK���n�<g��<�1�B$x �Abh#6M��1�=ާ�?�/l�?�4�!/|@��=s���gj�}�GТɳ$�"!��M�g�����s�WAX��n��	� �}�����x��.��W�l�2᮷���L��Hͼxi�&��{)���n�L$�\R�N8����ؔ����Ua�Li&��~�%)Z��4A!�뉅t0��yK$�JD�[5�u
�D�TG ]�$�>$�������J4Rp�<i���׷��d�f�Y]�_�*h s�@p�\q{�f�UZr���x��,�)Q��(tP�l�i����x�X��NinBi0�,Er@������LJ��$�Zc��+�-��&�m1A��|}~��a���}�rd��>,�lr�9A�
>�Rƚw�. �>�,��:L)s�",�K���d9�� ሏ�%<���du��9�IE�e�Gi�{4�G����ٺ���HL��K��O�NZi��F�X���s|a�8�Sqq�mT��P�':���������t&s�D�>�Tq秢���v̙�*xCaäY�N4!�z�K#��Q�.��y�ꬥOX����p�4@�
�&�Ӛm�f\�xӺ����������s�:Ϫ9=���2kzޙ־V�����N��w>����`���>��AH��%��(�E$"��RYh�y��K���H�M�a6�J��VI�ngɄ��>���|If9b"C�y�Ye���	���r���2d�$���Q��%�A��e��G����>����{����L$�C	1�ABh#O���9�9D�"�s�,���AW�$2L2,{(��N]�&Gm>(�HP��ҳ�4���0��x,�I� ��"� �h��3�4s��O}�劣��3*Y�L̓A�|�(��	!� ��'3AF���n�0�L4	ϓh9��,Er@�G��h�U���AZI�e��g(C������f(-q�}��sgʩ��f@����a�ziKx��(F�Qs���zV,��8C$4�I�Ib7�,�4�O��'�6������B���S���fN�f��5�ZG��7��di�B͟�>����e'/U륞ʫN�^�B��X�A|�,pa��=�W���'W�p��Yۚ�l�3om�wUJ��l����I�1f���^@݋#+ȟx�^>H"	��Zm��D�D$����'�d���EbE ��D2u"Κ�/+,�.���M~�A ��? �IG�YnQ�V�G���Ğ7�[���X�y�$�I�ir�9��s�z��D$#>� �2�+g�n��F]׹B��F�Y�V@@��4�>���G����Զ i>$�-����u�\��Rdl�Đ}�:�:ň�
,�͵0H�qG�5�*8�����x��(y"�.O�s�9D�"�p�8l/�o�>xQ���0���rdvÊ<)
ᆐo$��;y��x����TA�&s�/���4��Ӻ�����٠�����	-�B�r�0�-73a�9~��>���j(�,Er��i9Z9���?.�7w�:ߦ4��I����� ��s�v�z6dֺ�s�ߓ����pα1��C�h�>L����A�$ha;���+޳z�����V�fV�85��wW�5�g� gL��U�D�)�WK��.ܝ�۽Y�UX����4�`U�7��Ű�) ,��x�	!��O�B���>$�'�q�40������ϙ4hBe�ɲ�0M��=B�PZ$��s�*~����m���-�K�A�(�*��%�hx��wӑs7ٜ$Q'�$F�r��QF��l�4x��0�*��B�>s��4�c�Ĝxs19�?��5XЙ[��8���	��d[���h���y*����!||���Q�#�pJ$sM$�y���nwD�y��E�Hs�9�YrǊ����#X,�}�91r����I�ژ$} ���,P&F�^}�m���d���s0sr��Dc��ĚBs��N���[k����L����k>(�(C�X�1a�B�ߴ��s*�^�l3�����-���#�� �+t㢶�)��A~�dY�ć���Yy���.��|�zݩ��ÄA��c�Rn��-�ATKj�Wi�tΔ�ڹ]nu:�)&;�e��:��M�
̗��:{�w����A�ZI��jqy��G͐���/N��.? @/Z|����B$�Fc�"�Q �"@�S��ȭΗ+�����7=\:���:C�^c�w����ſ�d���G��nR(�ƒpf�D�}S^�!2L��k�r/���-4��zK9�������b����d!�� z��&����-��7�egzb�z/�&I��k,�Ρ}�D��A���҆*��H��		��5��v���B Dq��#��=�������BRK-A��sK����0��k�[�1�~�}��|˻�o(>*SH�8AY'�f'-4�i�1�si�����d�I ��b"DC�S���P��q}�~���L�	�<QdH�d���K<���x�����%�c�I�&�>t��簲�*�#�X�i$��wD�4l�{�|Ԣ���i� �b N�ӄ���٧N���5�~*1s��Zȯ��h0��	��`XC�YF*[�#̨j�vT���qvT���H����.�7Vsٮ	[4�w�6���Z�CnꈗzR�V��,�G�x���y���).m���-���'���(��	4���-U:V��;�k�$�Z�L ����t�(߉e=�����K�s���`�b��	�<Q����Ǥ��h����	3iA�.�	"�8��Zrt13}�+;~��=��g0��m0��!B4��O�����o0}�~��I�w{���$� �3�`��K-�Eq�&5p�M��芨�
L�G<a�'�r�H9��X��Qw�lϺ*{2����$�$�6H�<d�I��ϋg(C���ƛG3gė�ޜ�{���`3�(<�(�(r�z	r1�9���L��fc֝����P�I��˝b��ﰥ꫿ǒ0s�����4��y�-�4�M#��h��{�*�ێ������A$�X��r�H�`��+�\j���������H�� qG��M~v(�D��x��Գi��z)ײ<�N�,�j���<KD��N ��/�NڝVX�IY��
����IU7z��=�]٢Mr�!=]���'q[�KI�N0xk@
 	��AO��@@D3�������Aݔ��$�ι��|:ө�ޒ�L����	d� ��IC�ܩP4��P%fiG��Uue�+�a�4r�! ����r�r�B��9��/��ԓ��p�=�Q#�a%�刈I�0�8c/�>�|r[�w<�]L��22K" �$�r��>#g���Rw��Z w4���@�4��c�dAG3���w�c�Ρ�H�8�֜���Ŵ�������m�^y��F��8�����Ӕz�`�;>8�Ύ'���l>0qzO�ri9F ơ��pʰWި�#$�zK5�M �Ǥ�#��� �#����7q�Y�G��G��P�a:�����ۅ��|V���\	i�r�\lk�I�M<O���+���K�-�;9>�R�ܘ���
���ğ�U�j���1�g�M�5��\���?mp,Z$���]n��1�r��y�쭮2�:i]���/6�4Kp���s�]��Q�6�g]w,Ȭ�Բ����.5^�o@��5���|��W��3����yH�X)�Z��]�b{���<�Xzķ9�.�ڷ���%�{��k�pj�31hA�=����5�҈����l�{\u��מ�_f���F�38��ʸ}�[>(��UW��twVW�h<�$+�w����*�&gc���޿V���.�؎Y\��o�����j����q/L��.޼�\���[�=bg�zOz�M�:��u�@п.K]��k�����$q�q�����=�y.�Ιlꭜx���x
n_����/��p�K�Z��}]���k�V�@�)t���Z9��)�
P��{����{S==�� ��"�b�6q��}s-��F�W��4}��)��������F1��R���*,Z9>��jdu��kO@��U�ۃ�GFv���;��%4��=\��U`��ܥ��Ć�X�.v[xi�`�y�	������P�U{��� �&�%&fI$�����D���0�߷F�m�˯}�%�$�Im�����om��I$����I.�w3��痙e�������$m��4}�ܹr俙$�m����I{{{�'��WR�$�I{�Ye�I$�I{m����<�>�롙��:4h��"H!$JCPK2�f)�����S�����mp�ʬK\��O���ܕJoO��!AQ֓�d���6�[�7#52����Ʈ��F��t�Uu��1
D�Ԭ�XX�P���jPtoF��/8��{]��s��[{SN���I(Rw��T�����9h[�p��]��a+�c��ew
m��7�e�S�尹i�Y�y獻�@�w-HԎ6�`SNC���Hnzx2x- ��}���^�L]���{Gk,����6TY�͙x���g�(�	A��TuN)��W����ȕص{�5&����-WjA�}�����+kfN{�f��n�q��ЃI(���J�����J:�V$�L�X#6fK�gI�tK#6���j�{uy�N�{��M�����:2���!��y����z�6{qv���۬�7Mpn��V�<�����g.]luѸ�9gH}(��;Mֱ/�qɵ՜m<��S}م>�:���.��e�;TB�R�������ZK���b����^UΛNܽ��9��tW&���g�e�[��Մ�U�ٹ�M�� �����0\t�s�T�)9��,'���9��u��ʈ�@:2�_��Xi�jܪ��RVG)3t_��D���ud����u�=j��ɩ0�w��B��i��*Z�7��B�LVa<ErÆ�i���AF�b�������k��yqQ�J��]q���^&I��YUW�T�]���wC]}$b��b����"y�%V���'ge�'7����w&�ܳ�&+S���e4pYM�,����㽭��$vD[�C
�V�eЧ��H�Mæ�vItV�n��&��΋;�<������B|�K�H��(n-������alU*�9;8*�T�����(��(e���N�i�����[�C�R�w_M�֮����2���,w��-3A���S�8*�^�v[j�9m��T�0S4XF]�[�y���d�vJj�3g)���ń@���2��=�P�`w��/V}��y�T\�J�q*��c�.G�w_V��"y.�RUl���s���Rz��YX�;��0nǸӒ?].);��6fN�r�B���E��d�	�m@/[�.E������{f������KCT.�Zt/��64�xL����"��n0����'v��)��,;y�`��qG�A�8@�N��0_э���clbm.ȷ�U�jV�HZ�`.m�Ά�䀪Ԑ�ph�yml��ǖ-ʦKuxVQ��$<�1F�i����� �/a�E�I�����@��*���PA�䅐�F$MH�̂�t�a!��!%���# ����U�����r�@� ��M�N\��i�I�c�O�/lD`A�9'IF9e�G�Zi�3q���[�=U��s�0��19i�sƔm��x� Ჭ�>���x����r�e��d�	� ����1���3�[in|���,����a�u�\��5�ћ7u�g���L��DH� �����`����3K���>���x�v�ᢁ2$���a�A�9�u��"�_�> ��Pm�&Go�<[IBf8��=1^���4�����˧( ��	9��p��^��[�̻�c�K�i�,�j���g׻p��#�sj,Y���G���D�3{Z�!N���":��W�P�{���<�{��7, �0�0��W���Ȕ��N]*�_�=	�;����O1�Qn �����Z#�4GvyW��6K���i��(]�B�� >mEx2^u	H��%���f	H^�&����0Ā��@�T$ڡ^Z�0%0��,�LRB���<Q9wM�L�o�9����(E�	r�`�N~ct�g/��0���M�z���pH9��"8Y��꯯dG�* �[�I����s׾��^Ww��[�x��,F���8�d��U�I/$��3�i2x�,�(�4�c��8�c���1�F'14�qeab#7�A���aNߵue��P�{G<|�d���@�[���$�{�D��(~i�9b"C�5Ͳ˒iA��Q�ۉ�*g��xD||I�a0H�A��@s1���M�>w�]��D�����<e�Ez�	"�p�ʽ_MsiS(�]p�c�gLz�*�і��R*����K��I�?Bω��T�1���c�x\� `����GRu{tp��Qh�FR�e�sr4s�3��tFQ�'��3F庈V|�Aw�k~@�0e�&;\V�ϡj��u��R�e�R BV�g��	Q
�4���A���T�mI@�Ex���:��$A��WЉ�C(�NL��a��� p�o�+<#*S���z�.�u&�<8��|[����^�
��̱9%kP����8�Ɇ9i��o�{����;G4�<"�d8��H*����-�᏾F�=�c��Mda�$}���s���by���^c��#�5� �(�ʤ����"I(�Ow?l�8��H(E��!�d3�a�p�י��tY3?4��9e�i�{ � ��3���ݛ�q�1�ɜr4��!v���h�3<}_{�tY�}�~�<����5�|`�?��Q#�i#��P��蚥}���?{+ﴒ--�4�O�OA�3�1|Ο�:��i}P��/P�=��R:f]9 � �� �0�� �F�8M��DV�]U1�Õ36�-қ��ړTV�T8�� ����Nt�h��>�2��y�}v��B�����E�a�Tl�eB'��^�+�A$E#j�;w1Qe[���P�q!IihݡF�D��Fʵ`�^�H�AY��ڃ�ǷW�Hӝ��᠎�H���0�Y�B�Ib8�<��D�d�s,���`�� ��@X�L�5�:~�s��w՜�>2
GǮ
( �,p� �'�Nh���3;�_j�'N���E�-���i&뗃�Ĝf��EL`�� D�BD�9�>-ʤ�i0�i�f�?Gɼ8;h�vI�9i���Y��'}��mvfW0�z�rEU)+>-����+��D�O�=�m<I�Б��	4��9B6	r3�����$�K�Ɣ��v����@� ��O�o�3��O���c��}̇0� (G�;�a�Q�,�"w����|���]�������S��8�@Z�h��dh!�kP�@�~~::����B,�B�k#ֆ� Ϫt�Cs��A������1>���,��\A�4cd���7���̚32�pT��˱��lR���C2cJ��n��0H� FQ�Q&v�	4Hq4�:�*l�V(O�Arh�!��E"�@'Q	H�LYT�,�M��2��? ��I�]v%+�����At�7V_�x�M#�p�> �Oa�Ri����
���A��!AUj-���-
�4c�8�ǭ����5��������Q#�|Ig9b9��������\��ޤ��le�I���d�"<i$s�gG������o#,�$} ì���&Fx�5�h��]����� �$�<I�	̴��a5�v����>�0�J8|A���/.��oC�f�ʊ��H��3ҡ�6L-ʤ�q5s�7�H�f�1�r�3���-4��zKB4
�-�)ml]�V�V8��>*����g(C����6��n�U�I��[�Nx���}�'�Ǎ�8C�9,C�j
�[�[����-�Y���$v�Ya� �?�Y�T�0LW3+��NV<����ӛ�w�Õ��z�F`�GbP��q'����a�(1V�n@��-�"PQB��͵�fOj�T� $Yu��M @�,��ESq�(�!I�0'F��i3�u)(Q ��wA�ZID� ��i%�01I�Zݔ�^�L"IIF�ta%�}D�����H9��r�z	r1�<�3}��L���������rP�|I�0�*x͜=^�N֌24rN����珤�\�ܣJ��?�/7��^c�gň$� �� �Ri�śa�fϾ�&:�g�!A��-ȯ�,&�q�u/T�UE`Ŕ<�A(�ώ$�X����tÝ5s�>o{�����57�%��A��Hw+����LL>�4"G�>�8�A�Ѩ�.
(����Q�'×��H�8�sm9$�x�Ki8*x����׷��DAd�n_�.��z�w߯o���2�n ̔ ;�ۤ�;��_Os~���dQ�a���/7ob!��ϰ{�ˢ��)@���P�I�O:�g:wUN�J�ޮw��mG���Z� =�I�gJ�w*�±Ժ۵�4�_u�][D�A�L؃�Q�D;(`9m��&����mk����d�$`Q�4rE�'b��I�Cn��̔�@��>}��n���[#7u%/�ע�W�=TUUp!5��qʓKr�9F ơ��8i����x�X�c�2i�A�:KB=�9#A�'��ʘ�����������l ��Б������?>����24XZ(`#�K�A�(�ʤ����ܸ�ș�0�� DIğ��d9�A�z꽳*I��<#�w���ܣ�Zi�K�8���NF�Uvs37���<A�9I�s�śab#8a�0��v�����\O�����l��7�xy����8�I�-q����!�$9����\���t�D��b�Qaɂ$D|a$;��!��e��9��o�N�q~%g�D�|�[ ^�P#�~�5�:�*�RS�F�K^L��X Uu�:�z�
Ğw���ݏ{���b �A8A�f���5]Uu }�u�+T�ɴwz7��f��6���x�$��c��^wCuX�H@�m��t�VZ��� ʫY�I�F
�U:lHg�j�3�N�Q�aW�0�&^�ӭ��8K`���F�10�vn��Y��6��3���mFpQAc�4YE{~���j3���!˴����X��2����13�0�$�L�/�˪ DD���V�9�a�����N�ә�� �F9_'(��5�9��9�
4��k�a�9ϓh9��,E�8��<U)4��y ���r3�!��A��P���	8�y���v�ꊞ�f�C��1� ��A#_A� � G��8������@�r
(��a�T��@P�����H��{���rN�r�94|XI48AA'��[���V>�c�3"�sSH�>���DFI�C�̳���olEa_;=m<���I[�l/O�Y}�c���L�N�UkH�wU�ma,��2��42�,A�Kw�Xc�,`��n������N4���Ǜo�:]7�f���%Yt�UԤ��]��2äޱs 7��p+۷�!V�������������f1��c�\[[4��L�v�S"ˎ	5M���Rr8c-Ԥ�t��Q�����J�/$���6ں̾�.��3Y�n�`K�"�A����%�=�x�ߝ�`�4q&h�xIa'��.
M�'0I��]3��"�a�I�iȾ��Ab5��<x�wF<L�0��ȂJ*����(��8I�������d�`b��!ͤ��g-���i&�7v�1Ǚ��iEh�D��$$L�.s�>-�b+���1w�}���ǾNa�dj�r�p�-4����M��d�����>(�(E�$"�*����[9a�}Y�)Q�"��Y'BF�$s�sX�����5���o�)� �|����b �Q�?Q9*����W�e{���� B9��"����_���|�}dy�ZC��o���9ѯ��mV�I�V��K�%;󃆍4ha����n�kc-��Xa|N�Um,��ܧ5"�6��p�DoR5Ε$�*c�ۛ�/��K��p��8�!�,�����!�׉e�C��k��B�b�k�m����*���E��k�Y-պ��9��<���yo��չg��,�y�m�����m[)^Nwû8��؈@	1I���Ͻ93~��1'�<#Mr���YBm��d�����pÈ����9?MG�q���??��L�c3ZoqG|XX���	=�,�*���k�Y��UU5��7��i �Ǒ��&G�H79���}��ދ�0�V��<IPe�&�A��e��&,o�|v9$"��dH�㬒��&F3^�y�j[ww��T�9ˢ��>��H�$�A�a�ݾ����DU�p��rϝ���m%�0�I=�^p�a�y)w��s�����3��q͓�ܪNQ�9��߯�O�k�<�8;#8j��~@P��h�1�M��+su4w���4�7�Eo�mS)ڴ�_uZ�{�,�#�'{ʏ���"�ڽ�,��I.�C&�W�2������V�ȍ�Ӗ�oc�ct߯�껤.�a�x�f6�\�+�`����n�w�3�R�U����)��Y�N<e�Gv�[�ӭ�W��a��.mޠ��Ŋv�t��a�j�F��ɕ���=+rD=���%�;.fs�����
cHp��:�=}����NIZ�8�v=+���#��Sy[}O-p��w�ӝ�}G�%܉s��	3��5V(����	Ȭ3n�}���VnW�&N�z+�}A�4'�C/�����h9T�o��:���.���Y�J�o��x�hR��Dj�E0Aj������{�2�}�=����ή����Q9��r�oڥ���ͣ�����u�1�iv��$ו+��r�	�΢�Q�D�nI�w�Ԓ}2�g��{O	��h�/�n<�-�+�=��3r�#r���!�U�s���'�g�e�A�g�3ub��|}E%u��,;`C�L�n
6rz��rM�+MGAq�\C���w�#w�F����f�F��n��3y�%3w�W��+r
-d�Gl�s�u���7�u�ĸѺ6����UU^���.g�����}��h�� �uӜ�����r�˗$�@�7Ç	;�h�s2��&d�A9$�I%˖�l�Km��d�Ie�������^^I$��I?=����$�\��Ym��/2�m�K{���$�Ie�m�I.��[m��$�I$�c��z�������\�9�?��w$�HL3L7K7{}~�!�K.��S;�\t"����v�o
��`ǔ���m���ʝ�%�y��������s_��^���+�i ����8ei�we��C;���Zn��.wzp�Bo�o�� ��.�q{}�5RV��]rL+U1�Y���q�H��6�̕&�O])Y4���k.t7-�>AH��1f��/��:��|;rY����l������¡QU���Y$괎q�X�7,�o�|��+��Ֆ�uiWRS
ڷ7觺�)�oY&���'_pY�1��K������7{�utU:㛸�K�	9��3!��h�>��]�T��ɹ{\��RaW]Ʋ�ݼ짦���5Yٗ���eC���z�ޭ��iKN�v3:�I��j��-�m�\kT����WS�ΡF�{m��ٵ�7�f�F���}��oXi�n��m�P�Q�η��,'x�ݹ��
U���w�q5+&rU�����8�0�T�vV�M���r̝[���y�V�[<Md~ؖ�6��5Sn���:��Tѽh*}{�ֻ�M�z���S�
�]kf�����7w)\,Y��pUau;�%�ɭ�!Вzf��+��ܴn��t���b�w�J���I�K��K�w~��y.s$CO�1�B[Je�W��K�}��3��p\��V�D���:o2�0�s��Vh�<:���^�QӢl���\�l�'9a�P'L���s���z��c�����+0rƑ8u�(�Wd:�p�f�e�MEfZf�o�v�YF��w�u�%�h�T�#]�]�Pb�b�e5;V����g
v~5գ(:١��)[y:d9L64�ۢ�mﰾ�A��N�*�!���yb��A$�H�Q�7���cV���{N���c7�Up���7\l�	[}�z�U5��(R9��*���F�@��Y&4]�����}C:���	�r?���tr��>����6n�D�I�H����b-��K�b'���4��Z�l�Os^`T���,>�%Ѫ7}w[K�a��<�b#�֞�l�mio�{�a���}*�erHg_֋��0h�R���Я Q�u�f�9�r�4O+�.�㘁�l![ĸ�3X��ʆȬ�2�(����!n�,�(�t���b�X�e"����'t]�Xၑ�E
�b��N^���s���ꫮat�䲜��Ӻ���Uq�Vv�Jm����-]u�-cf�{���%v�=��:G��� (�w9���{���X�=Y�܍L�@�B�� E#�1/}�]��[�Վ�9����p�.��z����̄B��d�-��� �4�>��]Ø�9��m��>�P!肅B2R0�m���Yޘ�����j8���#1Tx�hr�lg^u#�Lck�|��%� ��>(��>���<���}h�[���]�&��=%��s��>�gޫ���/[�0��pp��O�$�NRi�M�d�]q��<"D$wAe�T�ń�g�$�;ν��b��Y���\#�|q�r�sH���K��7ԓ�Qe��.
M���H�
_���<��I�|,D	?�K8�A��r9��}�EUc���cl  {le� �߿f�E�]����n������ę�ya,�b�:����>@��$��~>Gܛ��sK�aw{h�գ�ۻ'w��a�<�1c�4��4pa�:IsvR�b����{r��d{��������TМ2�Ojԗ�{�R��$��[����@���a�x>L�!~����i �L���}Լ��e޺�ɢ����|��D�|�E2�d�M����q��5��}�������Xc} ���9x9t���N��/�&U=W�q	�Ԏ9�inU'(��j�&����S�1L�<a�g���H9��X���W׿J�z���ed9��
�%#�h(C���&�G�g�ޜ�W�h���H9DC�#�LA�Q�p�Ǐ�8�e�<[��PzKAĜQ�c�:�%p��7�j�xFU�&��$�E�r���I����o���Fb�o<K�I��n')4�i��e�s6z��h��X���YnU9ń�b M�Y�,�s�RNC�<G��s� ��	!�$�<��ǘ2����{�;N�De,]h����t�������Eyt9f�s��*:%j��M�y�c�81�rZ�,L阙���/��We�W�$eu�]�p�\�Ve�!�c����Grk���FyN���!,����֔^A�m�U6�Yu�a�w����.��k䌤1��yH��������� ��( �,D��d�rHE`�1�;_}�R��U^,�;�8� ��j0�.�9��/O:�|0�Ρ�H�>(��ӒK��8�����_�;�f�U� �K�����"Q!�\��ݝ҉����&��9�>-ʤ�x��l�����ws���A�>��P��G���]}�.����8������P�aĞ:�����ۅ�������"A� �Eȉ�(�(�m4��r}�U������X�8����d9���i�-[_�$�F"�9T|XHX(���[Q��O����_u��� ��{�Y�PE͓W��N� �L�8C,%o_xc�����-ΰ��0��a�|١-$�v���WÔ��+���'1�\��W:yl���f�h�Mܭ闚�R�J9P��2�h��-�P�F4�X�T�D/<̜}Y��(���!��JYAU ρ�,0��E��K�'h�!��;9�M��"#8c*��������i#�(�*���\�&��4q���7�"ٴ�>��,��r�<$�0���.���͛���3��l, �4D��$�rHE`�x���j�moۧ�}�w�S�h�8�AfQ�0�.� ��>��G�EJ�G��(��NI.�x���I{���\W�Xi�ĝ�^�]Q ��	?��9��6�>ߺ/���.���"��Y��8;`�ě����=���g����|d�"�}�9"�*���x�����>0�s�M�Ĝz���PH9�GO_���̺ꏐ��f�.o����Ԭ���\48�eY#aVG�oQyC�;2���^�k�Us��� ��x`�� X̫�����0��V��R\�d��C��V���M���Q�M�僅�� �t�!��k�"��V��x�D!H/",�y�b0@�4�^ڸ!DB��$VP�oh`�ǿ��I�#��E���b?���W���d��A�,F��K!�6�(Ls�ׯ$�)����Q��NUXI48A ����
��6�<���H��t�X�!A&�`��,ϧo�����ȸ�i�\�&��<8�anD�s1�]�}
�`I�u�h����Ğ��\��6Nf����L�����2O�$�WÒI�d#�o�����s��}w�&G�����x�.� ��G���zQ3� �/�K��qm%�0�ě�VxFT��g#�9wD����3���I�n<�l\����9��zv��ڭ}���$����E�V�m��D|��H>�쇧����|eZ��*�����1�0���Dl:ŋ��1cޱ�\i���������5����f
��Z*�؜�Νy��Ay}:� ������aK�,&��f��,���>��1��
���,��PPG�����W%�Z�IG��8;xsI=�Ri?3����=osy���x���H�yiT��il�36�@���q&BGت	8��8k�i�[��uD���ʢ�E;|x��,AsĖI����}q"$�*Y|z�(Lz#	=G3}��L�E�3�'���e��C��G��19�iwf�z�#�r.M,p���$��r�H,�Z��~��[�#���"��F��
Br$q�4��s�{o}��SW�6x�RC�Ip|�.��( �,F���}�$�c��I��O�8��X��������{�ߦ��~N����6Q��H��p!���<R�N���aȽ���U�V}�nY���Uku
��g�`��D8X퉴@��0X���[j�yһc\M:.��V�&�Jԡ�"�R�)�h�-���_j]�g"���>�ڂ�ۯ
1"O/:@\B����M$E��B(�|�T���,���gn��� _�"��@P��0^���!�fߑ�_tk�ED�Ԝ�ݨ�Ŵ� p�H$݂�s�$���Њ�½D�<HH��p㞓�ܪNQƐp��ŚO����I�^�&�sOIg0a'�ݭ�j����"EU)+���P��}�Ȉ�����A��Бت	4��8Q"$s9����I1����n'l,��(AqG�k��ߺ�����ӏ$9��	��B0�h�.Ӝ��q_{r��ϋ4D���> ��1ʑ��l����}
�͐xp�#H$���r��,%�<�_dN�j�n�� �b��/ �0�A��4��HD_�s�J"�K��RZ�<���{n�%, �0ǅ��#k�&s*��N�_'e�9��u�y�Ԓ9�  �U,6����:(��1�棻�j�:MR{R�7U�F̤(��= �>����B��D��� a��P�/��yXA�*�uU߅��2��-p�����Y�{_�����RHsI6E�P�PA�X�ɣ�G�s��L��t9�a�Abg#<u���d�O��g9�h9X�$d�(��NI.��*���ԗfg��X� p��	7�^UQ �fh}���yQR���g�C�l�[�I�0�j�o���I��lk�̃�2
M ���P�5��E78��}����`��R��sų�!��q'����O��wz.'��E-�Aψ=C�"=" s(��Ᏺ���"���Ğ��Ağp�1�)U>�<^�2�9�3�4�mB.�1:��� 3o��BW"�Z�+�f�X�G�ĚHI�VcGr,h�7�����|�#����9��7�eu^1������U�f+n��"��r���aƖ�)g��(� Y�&M���N[�ݎ���٫ծ��֮�D����ur�����o�&2#ğQ��NUY"'�(��}�z^c�g1b	2�*��H��6L,s�}�}�Lu\�����Q�YnU|Aa.X�q�w��RuU��8�i�D�9������N����r��z���>ϳ�EzJ.K" �<9$"�s�;������|i}�&q20�M�Q�9TQ�����11×��H�8�sm9$�x�Ki9���O���^��u�$AŐIW�r����Ჸ���ͪ*���Bk���'�Rr�<A�C��i���ǉ����>��H9�Ib(D��(r���}��MOI՟D���Ո)�ܤ׏���|�-�������2X�F���J�K��	>,x1h���1�0`��Aa��o_MerƟ�Y.�\�+n�f�f�ܐΡ[j;ͺ��̺����Qs~ŕ��G�� G��y��^�4A#շ_9��\��z��s����c�9�^Q�)�v~��v�+B/�P!�!����������ӇF��'��M�P�����T��Ҏ`=�N�A뙏5�� ����G��(1�ۜ�%%���G��v��<Y"&�f>�����dm�Wg3|\�}���Lr�vs��Ʌ���?�{8����Ɵ9U���b M���8�s�H�Ȉ��O99�vX����sȢ����>���#{JME�&�\�I��M ��5F�����>��_}�8�3���mF�Q@�c�sY^�AW�G��,q�NI.�|SABῐ�3 �cf��`�?���6cKlc�0f3նl��׮���l3�s��0ߓl`�����l����l���6m�������ٶ��;�_��_��z���1�
��+�)�@�fZa[mL(4��"�&֘A1al�X��m����̄رabhB�,[BX��i��FՊƖ51[5
�b�bB��+���b[Vf�(ZĄ�X�&%��b�(+b�-����[X��-��ZŖ"ňB,Yb�e��bе�X�E��[X�2hE��!mmbe�,X�5�����4�lX�!al�6�1bŶ!6�̱3!c,Y�e�����,жB2��be��,�b�Ѕ��X��-bЉ�ŬHK�B,ZĘ��ı%�X�"�X�X�"�BhYb��LZlհ�Z�bX�m	2k�Ak�b�akı�-X��BB�X�$ŬE�,D&��,�"!-�YbB�-�BŴ,X���L�f�#i���cX�,FX���F�k�k�kd�mbŉ��e��6���[Sm-����+*�Z��$T�J�iR�URT�V��YEՒ)Z�5m[)�3J�mM�6��j���ĶVj
�lVV)[jژ�����b��Vm,VձE2�¶��X�ն��6SaY�fV�-�L��6�e6���[51#V�X�Vjj��եB�Z�IZZ�*�Y�Ք�YESef����(���Z�V�D�mMMY���*[J�թ�l��(��JU�H�UQ��jԦ��J��j�QEe%j+jڍCSi�efV�V٫mM�j
�I��V��J$��SS+S*���QTՒR�����Յl+�H)��2���2XVaia����mmae�h!ab�X����e���L���aa���[i�mal��XBmf����L[�f-���6X[fX[1��FX[kV�XK

����2��Մ�A���KcMah#[kk	��0�k	��m[6�akmlAfk6�f�� ��VVm�K
°�����[XDXMae��a,k	��� �d�k	���a6���XXXXXBmb�i�XX�kmb��a5����2�F��L[-�������Ŷ�,XMal���h����XBm�a ���	�-a,"����	����X[kme� �a����������k	��d��ab��,&�Y�,LMaAma[j�XH(��4�AL+
mXVƓjbXH� S`�+
`���ia,-ak&�Ņ��mal���X[LKA,-`V
�-��ւk����a���e��m1a1�,e�����m�2�6�Afذ��[k6kf& �X�	���acA5���Ņ�md����b����XKi����5�h,[kd� �XZ�F����Kmm�XD�&-akm �,����k,-ak
� �+ �a�k	���"bm��,��4k	�XY���XX�m1lM��1ack�X[#kmm��afXFAl�Ѧ-�h&�-�XE���XZ�ZXS���Ak
°���XZaH+���m�	ah-�+mk	1h%������
�Y�XY�--��-�#XA���5��a�B�[i�k	��k	�ml��lX@������4�kf��-�aX[a6����Lذ�̰�k	�A3Le���m�dm�5��amaf���M1l�kXB�X��������-a�M�����"-�����A�XZ
�,%��"����E��a5��֘KXSi0�a&�K	����-����ڰ�+

�Z���,!�L�be����XZ
���[
�����6����w��6m��������6m����6��6m����6m����3 ����}9I 3� �FͰ?z߼�>��ٶ���`�#�����/�p0��R?X���A�l��!�l?�����1AY&SY��Ś c�߀pY��?�ݰ?���`I�J�HB�ZR�� �(*�[�҂J��%��˨  ���P@0��٥�Ê�J*������^R�ꪢ���{��*����� :J	�F��Ğ�T5����X����n��k��3��ioF��w8�Tx      i�JR���� 0L# �M S�0�� CF@di��h�昙2h�`��` ���S�MR�5Ta0��12i���i� ���       !Ijdȉ�����i���zi;�y�q�I���"�~����������a_�C�`�
Z��������������V��M�@���*�
�a(�2d*
��<~9�<������k�#P�kg����$��~����c�՗ �>�aRT��w����W�/���N�ʽ�&�,��ۓ2�d�t1�f\��Rݳ��M������6�wm�W��CŴ�ST(K���5�k�I�tۡFL2Sź�U}T�Ynސ��M���Ŏ�]��{3wK���}U^������_Rtu�Kt��Y��f�KO/b�a(U��a�>��ڗ�}F�Ӿ�خ�ay�ū3�Ke<�Sbs��6m�R�ڽ�aR��襰g���yݬJ�^�f퐝	*��-�/+�&L��m�u[В�J����p���h`����s�*s��1V������&ҙ���u�dX�-�hMV
e!y$Cs�_C ٖ��H�.eXu-�aԼ���OV��an)5����}��O��sկZۢ�۝�݀�Z0�$,�`����!8����y�<�/�<+Ѽ�N-:�u��_�T��ݘ�kYZ��\f��6=1���
f�f�A�8t�U��9HAD]F�j4o_nP6�]�.S\��У(�l�5ޞ����l��
��}C�yx]�Z�$��V�6�?wJޯW��w�I�QyOgӐ����=�%(H�À�	�.t{J��c!��4���C�Z�����fԬ��ʶٙ�e`��/$�|.%S�Z���� EɺV԰qS8*쪓߱,IR���350��knOk�L�-�d�9�0`�r�g�A��)��5W��L��S�wD�[.�UYq*#F�ԥ�������xĻ/|+�sjU���uڿ���xݙ�j̈Y9�Ƈ���QA	�{��쭥�N�N�~t�~�����i��!1U�"�S��{��)�9n��D��?J>����8.GG�@��h�9��
��:�u��������}�    ��� 
����������            ������   {������ �   m�             ���          ���   _wp                  ��              }�� ��f�.MF�)�p���zsqJ%!P��l*7B�Q�Pc�佾�Rw��=&n+�.�;�ww[ȌM�}�u��n�w.H٭��c�s+k%'H'/Rƽ���b�?{ӟ�HҺ�z��]���?V�n?u�ɳ�$��]�ce�WR��'��٨5\��nm�������|7SMe_��ۗ�]�(�S�:7,���y���a�v�tY����J,�td��ݾ��^��qe'�I��N�}��|�g���l\�]�?v�x��S�e�\��n�7	����$�4d�����Z����0�mk��4x��K��6��k,��d;[V����g'^cOz�r�gN���ݹڂ��優Ӛ����de�].���
�qA�1���S�	}ծҋ���W�̲�˹��Rz5X�d�[��˱S<%Gֽ-�M;{rם�+����]�/aǥ_��ܖ>��:��NL��7ջD�z0L*�k����F�{&xn���U�>��Kn��;����|�}W��Yhy-PLY���s�`�>�D��	��%v�I�pP��::�9���=��V{��YoM�<�j+ W5i\�B�4}��e{f�s3�v�r���q�W����'�¨��y}�C2!�83Ys�����|�t��{i�wu;�ܝ\�k�qF���Q�O�����զu�ϼ�U��z�V�v�v�T�����J��W݇��%��(��iY@ʖ6�U����*�A��;��3
'�Z�z��K���[�����S�
q��k[�CA,'}Oh�˸ؠ�5E���B�tG5ߧwuW�[��NۿK�ª������y�TA�]·����xu;����&�.��^�y���#�d.�#�-[��zN���(DZ7%i���*"�WtS���mU�w�u^D�Э�_�Q�O�馶�[5�.�r{ފ�_i�V{V�X��A�A) ��r�y��G)�k8���2�:������Ƭ���30���{9嗭G-�}x���J���M������@9�W�o�pe��V_�*M.������4�q酕O�Y�j9��;i.�S}u���� ��e�u샸8ݽ�E��頮�:��w�m����kz@����hV;v_��y��ehWu�@������۾�|���_�t���]����kd[;VQ9[Z4���=��|�
����N�Rc""+c��v��2�P�D̘Z^��
�I��^�8g���?�Ҧ�Q>�v�ʚ������XU�I+�i�^:{�lC�[e�����}�=yq�J�B�nde[��bmk�`Qt�_pe��ù��.��R]��{����n�7^�J7_�`�ǹ�Ϗ���'h۳kQ~�~���}'T;�%�ʽ���H����շO���2eܕη]�˫G��������YX�޴��1��2��t:�I�8`��X��-|:����p���d�GUݙZ�^��2����{�&�� ��_D�{�5��+yVf��Kb!R�����[g��p���o3���2^Awյ)֝M�ߟA]�V�<�:Q�c���Lr祬]��}|k澙5���ݸ���v;q��Ҧ�K���*�k9BwS��1h�s{H�x��w�� f�����>	�HM�b>"����O�?���  �@  	D	B��"4�u������ޯ���9x�N����:�_Y�y�z�f�y�v���M���e�۹�w s32::�|[x��q��`�� �v����HUm���u�q�OGH�Xh�"����f.FU�Y4���@za��G�#�yZ@S���Uo��o�Y�(����E��󍴛�Daۉ6�F�:��� ��c������'���@�uΞzx-k<oe���X�ھ:1 N��E�Y����\�˒�қ;����{�b���)�4њz���M�x�v-M`��p�˓�
����N.W�^ͪ��zҎ>�3�=>�̶@Ȭ���52���m,��+^����?f�>�v��۳� ���K(��+�7d=ĉIǍ݆X(0q�ż��7ey�`ʡ�k��3^FT(7̛�s��]X��f�a��	 ��]X�	IꮖNQQn�i�P�%U�o	�oS�	���JK4ogl��� �bQd�M�7�gw&[��~/�mzw5�*R� f�v:�5f�V	ac��\x��v�y�:Y���{���"<`�ye\�q�,��QB�txekS5�Ψ������K�^5�BH@;���/fz|q�Z\�3P���&}z5�%�ΜJJ�P�o�P%>C��'<Y�u� ������������]>z��N�*� B �T6����K�2#K4e%�Ǎ�ו�Pxk�J���ʸ�]籬U��ev����T]:V%C�$��>���z|u�m�-B�rˈ4Y7�L����T`���%ℱ=B�Ĥ���X(�@2����8�ۛ��^w\*�e��%P��?�f3����g�B�!�\n>���O�hZ�b<��mOu�3R}[gr�t��vDL^�
��:1=~�<jH�=~����q�����/��f�W.���17�؅2 6��w  R�`�4�LF��`y7m���8�����R5�0/"�C�]+���f[Ժv�8.fc�x��-���V'9�ʸ�}:�nɞ��}/ޯ\*$��xOʆPE�H�H�(㳍n��@�%EK}��Q;��ϛ���笱+аe�jx�3��˷�.��?%�!�Bk1z�Hsd%C�:@�Q�&@���))iF���8�t�%���!(JJJ�zi^�.Hu���(�$�&O��^v����)���=%��z������9���2`0�f����'��:n!^o{T��[�����:�nДw���R�*�4�>q�A��]�S~u��]�;ơ9�R��(��j�#m)��%	@oVBPv�#��^��t��J�Ր���K :q׮��%	GH���;Ò�%c�@�ĕK�L���H�4:�J�&�K��S���(%(�H�Gm��wpA� �(4��)J �dJ��҆����(J�,�@Y�I��{�|�{y�$2Zg�j��(�$�&OX�����!)l���<ˑ�	I�:444X�z��,��(J9��m-�2

��8�{@e߷m��!(���%	[�u��Hj�J���;��J5�S�r��7�!(:C��#���Nt�BRRw����Ր�%6�iu��9'YrJ��5dq�}���!(�!(JJSn��������̿��=��G QX,��(J6��K��ݴo	BR�	BZ�r9����2���vZ���b��_"+���z3�f�G缸q7�|(�����[��]x��N��m:ͯ��?gG�ug=eg����,wI02``��Z��;9 � �����,�Ǳ��Yݗ8�_;�
��N���d��AA���0s�&w�2��(Z^3�`L�# �J����ۯ=w� �
v�E��.�90�N9�6!���;��Ӎ���`�����|�AMVϪ%�	OŶ����D҅F�%���`�D<_CH���,�єRO,��-��	}��	Y������C�s}9}]O��%��,(���`5�,*f7�0�r$X��=	O'n�Y�>0Jĺ�e+�׮��`��ݔ��ዘH���=����>>�	{u;0��7� 2���q�X��ױ&_.���%������x�:�vfM#*.��I$�K�T*�ffA	oV���FʇI�Gf��u;ig�������L�A��yЉ�N'�تQ�o4d��*�\%�y,�8�h	[�d��ħ�L���g4��R'vd0�d�G���+�937��N j���2�A��s�/��k͹�φNc�X�MyN	@�楓����Yb��G:���D�W��������;��=�2�^�fh�)n�<i���֯�x���Iu��7{Q*]��ܳ������iV�Ш�I�T��F���[iW>���һ��-0�x��Y� H  #���#U)�Tv�f������׾���g\��W㫯�y-|�u�#�O|��K�ս�Mu�Zj�i!�	 ʗ��l��->��|��$߆���۲�_�D���|2����z�!��tH\+5�X���Ȝ�닊���/���&���|��y�o:j�V�(i��(��*$ѓ�0�LcЬBHE�� a�*�$t��:�{U.x��G����d̵�);����ssPxl��\C.���uӌ����0J��k��͏��E�{����(I�q���Vgz�'u͇��E�.��0�!K�(K���V|N�2����8�/.p���T:YoU۾�ksS�H@��f��~�ޙW��B���p,�C\����+tѯ�^:�pʊ�&�%Z�gd��B�a��O/&)AQ�$�->_*���?ٕ�'UA�:N�-�a٬鼨�
��k:xJEE�ľW�'�O�/~���|�&���~q��l�MB�Y��������wr�]V>2�W1$��w�p�M��J����,0����J%�Ly]z|(#]�s���`	���3���������1/��lS�}y��?��T]�xIi%+�q7*�5��ӉX�d��� I�Q�4��`��);��Wz�(���JǌX2>�:��vn,R�@�at/�d��K���+>�K�K���Ň-x��XVŠ �)�5ĺ��v�.0Y�\�#��k.f���FP8�	Gξ`�
뼖����7\Q��t��+��|��߾��_�?U���h�Y�t��(0N3UWO2�������^�q�¯rR��]s��5ۥ����2�u��xT�B��v���E'ف��1�<�01g��������&n�{
�������ؼ��U��~Π��B�zym���Y��	��9z��\�"<#���nz*N!���w�� �e�_�8 ٙ�� TE8}"^�y��]K̚z��,�I][\to
���\��@⚶-޸�Τ�N�ތ\8wM����[����M�O�x�K��-^, �r	gIHO'-���[ؚ��\�I��4�N�������i�S���s��񁽨@��nwDa;Ö�T�|vg:I�l����άњj�|/2�z8J��6a��6�嗄�SX�)�^<)�9�� z�n�iw�ڃ�mMV̢�TLY�ˏ��U�gyմ��[�Ic(�����M����R�t�7��%��Ms������-\��}N�=����ݣ�Hl����}If�_Qz���\�'l��+
p�U�\U��R��L|1Z[ѣ��u6%h�`��$|�ѳ|���9����#�v��v�3z��`/<$�WEJ�Nޙ�Ö�+�H)�6&�yn�����I<�P�UV�������g�u'��2�wX9_4�j�� ��M��n4d�׳Y�ݜʹ�y{�������=[��qk��N�.�i�o?)nEi�^k���W�V�M��ʓw��u;�܎���Y������l��;:~8ox�J�ڞ0�U�UUW�����	���拏�wu^�"�pg�|��°�ه}��1罷����VV�DA���b��ο*�SX-f�w�_��yEO"@��.0���c'�r<©Z璙̏���8��!#!K�?3>PH�c�k��:�ˌ�[����I6+�t�Y5��t[�}~�D�\�M~~����'�Ҧq=��?o?k��nC�n���;f�U�ȷ�Ծ��      !h�8Ȓu)�J�d[���Y�1z{�����N0~�孎��mup���з�'��Ur���$�0��{��}�{w�~?�Kԗ�L�:Gh(v��㦃'W������eT�L�P�5)�C&*a��Yj-dH-���ِH>��{p�r�:��W�)ʩR͔�V�xWe�a��@ܼ�kE��0jڅ������i����߀�S��������m�d�r�+I��P�xcG�z�rR�<~���ﾣ��z���ݔ��.m�D���\H���q���\X9�[���y�ѯ����Ѭ��{�w&˕�־��[�R��䍷�=H�h�~hL������S�)����oڕ%��yy�jzYQ�tg&i�����J������n��i��gYx0�u�W�1G��g����}�羗~3�j��Ye��>��?U��r�&���[_��x����s�����՛�����qP��`5'������>�=��U%�ff}�y�����_�̀��������� �����.fq-�V�z��꩔�Trg�s��O]ϙ�۶��{�Wd�a5qx��c��30erjH������	�o�kT���rx�l�D �j��T��������z e�̦n�����i�*ݛP��U #h\��ETƳaBS�jFh���A�^�-��Y��U3n�m��ͻ,�/2�+&�^���@\v������s������8q8�i"x:Z�.�`�Ii?�ɷ琴�Z3}����{Cw�ʹ�XS�G�=�Vu��+PF��}`��̦o���w\n��:������������  �3;� &�G����TR���]3A�����n�y�Xu�y����Ô�hw�xL�d��*)�ׇv%ճ���7��Ӻ���R�Y���uc�<.C�Q*����"*�9��%�	��@�"aA���!ݡ��N��M"h{yB���>)�P}�'���1��Cy��F'�#4��ь����Y�Os��z3��0�\wʳ�|J�WD�w�����=��^� ��}�ص�{�y3�+�����UY�ɷ�o�^�;KE�X��1V���k�)͡����K�M�Ao �����X�%��yPq6k�P&3b���N��G��:�Nk�9�O�=�8�0�u���}_F��V��ׅ�TdP@�7J2hOUp��m�)�I��ej�*ɳ/x��l����+,�=�޺���:�5���ُ�i6���}��a⯳7�/aY�y*�B�}Ʌ#�k&��]݆�����i��7�v��'�"鵍�f�y~+|�ճV�>S�����kċ�1��|�;+��i���=��:����͂�,oߐ�^��ܜ���'UU�o�A���������kq!||1�:��l�u}�ܭSM�	���߃5�����!�3����쇨�6H���4Ԓ�K��O��\\�J�m ���X�3r���(��Qr:$�=�^~�)���fM.��<���{�����;ޙגv�L��#j�g%D�v3�K������O m���̲����	��}ٔ�� $�  7D#l����	��W3�+n�)������XQ���{�3�u�W��c�~}�2��Č��I
�!C���o�����Dʝo?����&��QU6%*�w$_%Wn(�ֿ�UBK�v�7N����U��N�V��};��i�����R�#�&o<��:�u�j�N^�|��M������},������u�6����%:����}X3lP$��*.�mQnb%ꖸI�����ս�˿ߥ�~�ٻi���1�!�y�gOH�a�V]�i����=)<�][���h��`^�o��\S<o��v�I۫��x����|{������:�H��2�*Γܶit�֏���7_T6�`����X��{�)B�r����1���2X��{!�J�DyF�)(�HUy�|���y)�yΪ�Xy�&4j�}�{����CL#��K����iW�Vo�����WE�-�����������u�&��>t��Fs/���q�p��Y�3�����U�u�w��zl������2�A��2�TJ)�ѿJܴV��Xve��͐�ox�E�����������;.N�	�D����y�}��yC{��*,�B�{�Z�.7�[��N�@dby�v�W}����&�Y�oRG�A�Ë�z�j�g�)����Q�td���=w���v�������.b�������f�WZ��Cc�ݏ������͗��LK&;� nG=K߯뛏=��v��[aA?_��`�T�r���y��� ��K��y�� m���  �D	8�!��`��n	]u���ͧ�N�]���J�XJ��Y"6����owJq��TJs�vndm��t[y�K:���?J;A/����J-j���l�e�j&���:#�X����/��[�x��T�&�����8M����NaG�j�g�, �i�a��p�����:'p�{jH��dj���������Ҷ���Ո��<�q�Q�n�<�g���U�(�̏��k�i2#V*��Rٞ�R[��W�t�v��$�����֘O��ӻݏ��@��K����R�����A�z�f'��j���x��SRH/*��3h���m�ɰ����VD���Ԓy�e�� x��q6�=o9�7���ʙ�J�O�Ҏ��>�w#��X����o}��|+�V�>��o�v�c+�����(�{�nE|�"ο?t�������Ȼ�ռ��%(aaB��ZEu��ߥd{��@[v�y��2�x�u����]?3��5՚�n����p !�q8�B��#B�Ve��J7+;r��R�k�4��f�њy�m�
��O~��3��v�T���̷d ��3C�&(X����}�2��K��d��G�yJ�El�<ۧ=�a�o]� 1>ٕy�]��c�ż�T d!0"�X*���*���� ��@v���}�d�����Ȧ�p{IiW�V-�w�t�T�;�ɾ�n��3y3�7���s�00�&���&"i ����h0�]�N\���2�s|��ޞ���|6�:����6J愯%���K���So�������vEJR�ZM��6=����<��\x�\˝D����L�h�����fB��N-�9wV˿Dbb���"ys�6r.m��Y?lz{{�� $�  F�&��%)P̝�]{{x�.�Z^��\�A%���m�� A�U�y:x�ZK��~��҈j�(e)���ޔW���7�����Wj?:j��)Su����Щۦ�үaT��r����Q4E�T�N��;�L4
D1�q�K�b��V�k5m;k�&���d��t��p}������ݔ�h Ʌ.�M4A#�&@ST9&M4�RT*�{`n{wޢ<�1_eO���sy�F��}Qpi���)KL��tg�/{�u���y��c�@�;�L �!��q�D���;����q�	�=�E��+��j��'q�{�I�M]�� ݷ��.���c���m�ɈU:I}M�r:�8��IQD�O�m*K�ԏ��no��?������}/nD���A��?:3ɰ�?:�	�UV���[��?w�һ!���M�I$�4:�(ڌ32�3V%��lfZ3,��Q5��
�Z5��Z��j�,p�ʊ�)���`�%��B�b"9�s�j�{x�IU�۲�%޲�	�U�3�n9/n����U��N;�BI�;��C�U=)���Z�Ɵ�R��@O�D�N�ɷMST�j�UO��ۏ)��m����kp�<����a�ϋm����+���^���Jv���-�Z��d�Uf9Z�Zk�QT�����n�������3����qm����Xͣ}��m����l��e�L�I�*yu�<���,i;�
m��ڒ��R�RQR���K�!�%I|�i��3};_��Y�&9o�g+�:L�y�|�)=����4z��<K��OI~������ߎ�~I?�$��Q�����-�R_�S��x�MB���bCr+�a�^���ӓҐ®'q���my��j�n��XvL�����h@C �ي4�W�I��˞Ė9�9@l����h�nX'����0e�{ì0��ɠ 1��y�fw�}�a�կ^�����Gm�7�f��F��bo><+���~��g�)\y����ʥړ^� ǕW���r�����z��|�A~s����W�p�j�����|�C����O�<o��Y��sm���/����;;޵R�=W�e��F�q�ox^���YA���w���� (o�3+6��� 6���  T2�"qL��&=��N��F�!BoX�}�N�3�]m�q�/����fv�{���y45��,���u$3#^µU�9���1�ϸ���fY�[�Y� P%�D	�R$�����fSm���uA|����_[t�E_(����qڟǎ�9���E/´���b�os5\6W#�ߗ8|�u.�L�T�Ȁ�7�v����h.��Tj?-ݜ�����+���#y�z�p��{IiWn_����4\X�=�����w ��
Υ�qj�v�f�k���O�\vQ0m���ڨCo�F<L�7�%��ﾪn�r�~�O��'6����d��f;��g$F���0"�g��R)�;�5X�kG��Z��Loy�,i�W����CX�~�C�Q��ܯ�߄�T'3�P;�-�C�������&莬�{�-?G�B�S�������(v}��xY�W�~|�s����������s+V"�r����jU�Vn��E��x��6͏�v�Q�y�����y �LӢ7	����H�b�����vU�{�~.��/tb�JǬKݝX ����vo�1�
Ǚ8��^�*aY��{ �R����0�\�U�f���f`7`��I�g�P`&�3l6ϵ�1�`������pJͨͷ��3m���~C/7�yߍݺMW��Ξ���1�ϟӻW:��~��$̗����~   ����,��!d�����f�c����A��re��6�H����)?,F:�j4y�ɣXqh36�����(�&��;�ޏ�AA����t��:�p�Hv�N�z���͍~x����|�{H8�尿���Ɇ�����8������l���/W�y��C��`/��좂���������v>�~b.���C�������� �����?(_��� �7=���t�z�q�7~�����_�> �������z�= ��4� ��᷈hƈ���q��w�Up�LQ(
Z "`!� &����@ZU�R�` 		Xe� &��Z �&U�(
"D���	�"�"Z`$ ! )e`$`$BT`$ �E  T��H	��Ia�� %`!�H
EZJ �E�)R��D�X�X���(��P�(��aD��]�O{�:84��� �����w�c�|p
O��C�8~���|����U�>c�>�����Ч��|P����ߴ���Q�(9˰X}{������? ���0]�~^ߠ����������������� �@������,�������=��� �}��C�e~�=��A����U_Vn��_ q z? �84+���/�C���y���:1|��� (��U��8��Wn �ӵ�l��ǌ��l��ra�{wU�z@�������C���~~'P�X���H� }G���^�x��� Y�N�@?Z�Oh�� >w��Q�����g�q�t>�����;���� ��>yS��������M��X}��ǈ�TA��T<<��7G����凇��~!�@���y���!�p���FA�$"{� >�8��������Sփ�g�����x~� �x��+�O Ϙ�U���{����"�(H%�� 